library ieee; use ieee.std_logic_1164.all;
use work.gumnut_defs.all;
package gasm_text is
  constant program : IMem_array := (
    0 => "111100000000100000",
    1 => "101000100011010001",
    2 => "100100100000000010",
    3 => "101001000011010010",
    4 => "100101000000000011",
    5 => "100001100100000000",
    6 => "111101000000010001",
    7 => "100001101000000000",
    8 => "111101000000010001",
    9 => "101000100011010011",
    10 => "100100100000000100",
    11 => "101001000011010100",
    12 => "100101000000000101",
    13 => "100001100100000000",
    14 => "111101000000010001",
    15 => "100001101000000000",
    16 => "111101000000010001",
    17 => "101010100000010001",
    18 => "001000010100000001",
    19 => "111110000011111101",
    20 => "101101100000010000",
    21 => "000011011100000001",
    22 => "101111000000010010",
    23 => "111111000000000000",
    24 => "111111000100000000",
    25 => "000000000000000000",
    26 => "000000000000000000",
    27 => "000000000000000000",
    28 => "000000000000000000",
    29 => "000000000000000000",
    30 => "000000000000000000",
    31 => "000000000000000000",
    32 => "111111001000000000",
    33 => "111101000000100011",
    34 => "111100000000100001",
    35 => "101010000000010100",
    36 => "011110110011111100",
    37 => "001000010100000001",
    38 => "111110000000000101",
    39 => "001000010100000010",
    40 => "111110000000001011",
    41 => "001000010100000011",
    42 => "111110000000010001",
    43 => "111100000001000100",
    44 => "000010100001000101",
    45 => "101011000000010001",
    46 => "001000001100000001",
    47 => "111110000011111101",
    48 => "101110100000010000",
    49 => "000011011100000001",
    50 => "101111000000010010",
    51 => "111111000000000000",
    52 => "000010100001000110",
    53 => "101011000000010001",
    54 => "001000001100000001",
    55 => "111110000011111101",
    56 => "101110100000010000",
    57 => "000011011100000001",
    58 => "101111000000010010",
    59 => "111111000000000000",
    60 => "000010100001000101",
    61 => "101011000000010001",
    62 => "001000001100000001",
    63 => "111110000011111101",
    64 => "101110100000010000",
    65 => "000011011100000001",
    66 => "101111000000010010",
    67 => "111111000000000000",
    68 => "000010100000000000",
    69 => "101011000000010001",
    70 => "001000011000000001",
    71 => "111110000011111101",
    72 => "101110100000010000",
    73 => "000010111100000001",
    74 => "101110100000010010",
    75 => "111111000000000000",
    76 => "000000000000000000",
    77 => "000000000000000000",
    78 => "000000000000000000",
    79 => "000000000000000000",
    80 => "000000000000000000",
    81 => "000000000000000000",
    82 => "000000000000000000",
    83 => "000000000000000000",
    84 => "000000000000000000",
    85 => "000000000000000000",
    86 => "000000000000000000",
    87 => "000000000000000000",
    88 => "000000000000000000",
    89 => "000000000000000000",
    90 => "000000000000000000",
    91 => "000000000000000000",
    92 => "000000000000000000",
    93 => "000000000000000000",
    94 => "000000000000000000",
    95 => "000000000000000000",
    96 => "000000000000000000",
    97 => "000000000000000000",
    98 => "000000000000000000",
    99 => "000000000000000000",
    100 => "000000000000000000",
    101 => "000000000000000000",
    102 => "000000000000000000",
    103 => "000000000000000000",
    104 => "000000000000000000",
    105 => "000000000000000000",
    106 => "000000000000000000",
    107 => "000000000000000000",
    108 => "000000000000000000",
    109 => "000000000000000000",
    110 => "000000000000000000",
    111 => "000000000000000000",
    112 => "000000000000000000",
    113 => "000000000000000000",
    114 => "000000000000000000",
    115 => "000000000000000000",
    116 => "000000000000000000",
    117 => "000000000000000000",
    118 => "000000000000000000",
    119 => "000000000000000000",
    120 => "000000000000000000",
    121 => "000000000000000000",
    122 => "000000000000000000",
    123 => "000000000000000000",
    124 => "000000000000000000",
    125 => "000000000000000000",
    126 => "000000000000000000",
    127 => "000000000000000000",
    128 => "000000000000000000",
    129 => "000000000000000000",
    130 => "000000000000000000",
    131 => "000000000000000000",
    132 => "000000000000000000",
    133 => "000000000000000000",
    134 => "000000000000000000",
    135 => "000000000000000000",
    136 => "000000000000000000",
    137 => "000000000000000000",
    138 => "000000000000000000",
    139 => "000000000000000000",
    140 => "000000000000000000",
    141 => "000000000000000000",
    142 => "000000000000000000",
    143 => "000000000000000000",
    144 => "000000000000000000",
    145 => "000000000000000000",
    146 => "000000000000000000",
    147 => "000000000000000000",
    148 => "000000000000000000",
    149 => "000000000000000000",
    150 => "000000000000000000",
    151 => "000000000000000000",
    152 => "000000000000000000",
    153 => "000000000000000000",
    154 => "000000000000000000",
    155 => "000000000000000000",
    156 => "000000000000000000",
    157 => "000000000000000000",
    158 => "000000000000000000",
    159 => "000000000000000000",
    160 => "000000000000000000",
    161 => "000000000000000000",
    162 => "000000000000000000",
    163 => "000000000000000000",
    164 => "000000000000000000",
    165 => "000000000000000000",
    166 => "000000000000000000",
    167 => "000000000000000000",
    168 => "000000000000000000",
    169 => "000000000000000000",
    170 => "000000000000000000",
    171 => "000000000000000000",
    172 => "000000000000000000",
    173 => "000000000000000000",
    174 => "000000000000000000",
    175 => "000000000000000000",
    176 => "000000000000000000",
    177 => "000000000000000000",
    178 => "000000000000000000",
    179 => "000000000000000000",
    180 => "000000000000000000",
    181 => "000000000000000000",
    182 => "000000000000000000",
    183 => "000000000000000000",
    184 => "000000000000000000",
    185 => "000000000000000000",
    186 => "000000000000000000",
    187 => "000000000000000000",
    188 => "000000000000000000",
    189 => "000000000000000000",
    190 => "000000000000000000",
    191 => "000000000000000000",
    192 => "000000000000000000",
    193 => "000000000000000000",
    194 => "000000000000000000",
    195 => "000000000000000000",
    196 => "000000000000000000",
    197 => "000000000000000000",
    198 => "000000000000000000",
    199 => "000000000000000000",
    200 => "000000000000000000",
    201 => "000000000000000000",
    202 => "000000000000000000",
    203 => "000000000000000000",
    204 => "000000000000000000",
    205 => "000000000000000000",
    206 => "000000000000000000",
    207 => "000000000000000000",
    208 => "000000000000000000",
    209 => "000000000000000000",
    210 => "000000000000000000",
    211 => "000000000000000000",
    212 => "000000000000000000",
    213 => "000000000000000000",
    214 => "000000000000000000",
    215 => "000000000000000000",
    216 => "000000000000000000",
    217 => "000000000000000000",
    218 => "000000000000000000",
    219 => "000000000000000000",
    220 => "000000000000000000",
    221 => "000000000000000000",
    222 => "000000000000000000",
    223 => "000000000000000000",
    224 => "000000000000000000",
    225 => "000000000000000000",
    226 => "000000000000000000",
    227 => "000000000000000000",
    228 => "000000000000000000",
    229 => "000000000000000000",
    230 => "000000000000000000",
    231 => "000000000000000000",
    232 => "000000000000000000",
    233 => "000000000000000000",
    234 => "000000000000000000",
    235 => "000000000000000000",
    236 => "000000000000000000",
    237 => "000000000000000000",
    238 => "000000000000000000",
    239 => "000000000000000000",
    240 => "000000000000000000",
    241 => "000000000000000000",
    242 => "000000000000000000",
    243 => "000000000000000000",
    244 => "000000000000000000",
    245 => "000000000000000000",
    246 => "000000000000000000",
    247 => "000000000000000000",
    248 => "000000000000000000",
    249 => "000000000000000000",
    250 => "000000000000000000",
    251 => "000000000000000000",
    252 => "000000000000000000",
    253 => "000000000000000000",
    254 => "000000000000000000",
    255 => "000000000000000000",
    256 => "000000000000000000",
    257 => "000000000000000000",
    258 => "000000000000000000",
    259 => "000000000000000000",
    260 => "000000000000000000",
    261 => "000000000000000000",
    262 => "000000000000000000",
    263 => "000000000000000000",
    264 => "000000000000000000",
    265 => "000000000000000000",
    266 => "000000000000000000",
    267 => "000000000000000000",
    268 => "000000000000000000",
    269 => "000000000000000000",
    270 => "000000000000000000",
    271 => "000000000000000000",
    272 => "000000000000000000",
    273 => "000000000000000000",
    274 => "000000000000000000",
    275 => "000000000000000000",
    276 => "000000000000000000",
    277 => "000000000000000000",
    278 => "000000000000000000",
    279 => "000000000000000000",
    280 => "000000000000000000",
    281 => "000000000000000000",
    282 => "000000000000000000",
    283 => "000000000000000000",
    284 => "000000000000000000",
    285 => "000000000000000000",
    286 => "000000000000000000",
    287 => "000000000000000000",
    288 => "000000000000000000",
    289 => "000000000000000000",
    290 => "000000000000000000",
    291 => "000000000000000000",
    292 => "000000000000000000",
    293 => "000000000000000000",
    294 => "000000000000000000",
    295 => "000000000000000000",
    296 => "000000000000000000",
    297 => "000000000000000000",
    298 => "000000000000000000",
    299 => "000000000000000000",
    300 => "000000000000000000",
    301 => "000000000000000000",
    302 => "000000000000000000",
    303 => "000000000000000000",
    304 => "000000000000000000",
    305 => "000000000000000000",
    306 => "000000000000000000",
    307 => "000000000000000000",
    308 => "000000000000000000",
    309 => "000000000000000000",
    310 => "000000000000000000",
    311 => "000000000000000000",
    312 => "000000000000000000",
    313 => "000000000000000000",
    314 => "000000000000000000",
    315 => "000000000000000000",
    316 => "000000000000000000",
    317 => "000000000000000000",
    318 => "000000000000000000",
    319 => "000000000000000000",
    320 => "000000000000000000",
    321 => "000000000000000000",
    322 => "000000000000000000",
    323 => "000000000000000000",
    324 => "000000000000000000",
    325 => "000000000000000000",
    326 => "000000000000000000",
    327 => "000000000000000000",
    328 => "000000000000000000",
    329 => "000000000000000000",
    330 => "000000000000000000",
    331 => "000000000000000000",
    332 => "000000000000000000",
    333 => "000000000000000000",
    334 => "000000000000000000",
    335 => "000000000000000000",
    336 => "000000000000000000",
    337 => "000000000000000000",
    338 => "000000000000000000",
    339 => "000000000000000000",
    340 => "000000000000000000",
    341 => "000000000000000000",
    342 => "000000000000000000",
    343 => "000000000000000000",
    344 => "000000000000000000",
    345 => "000000000000000000",
    346 => "000000000000000000",
    347 => "000000000000000000",
    348 => "000000000000000000",
    349 => "000000000000000000",
    350 => "000000000000000000",
    351 => "000000000000000000",
    352 => "000000000000000000",
    353 => "000000000000000000",
    354 => "000000000000000000",
    355 => "000000000000000000",
    356 => "000000000000000000",
    357 => "000000000000000000",
    358 => "000000000000000000",
    359 => "000000000000000000",
    360 => "000000000000000000",
    361 => "000000000000000000",
    362 => "000000000000000000",
    363 => "000000000000000000",
    364 => "000000000000000000",
    365 => "000000000000000000",
    366 => "000000000000000000",
    367 => "000000000000000000",
    368 => "000000000000000000",
    369 => "000000000000000000",
    370 => "000000000000000000",
    371 => "000000000000000000",
    372 => "000000000000000000",
    373 => "000000000000000000",
    374 => "000000000000000000",
    375 => "000000000000000000",
    376 => "000000000000000000",
    377 => "000000000000000000",
    378 => "000000000000000000",
    379 => "000000000000000000",
    380 => "000000000000000000",
    381 => "000000000000000000",
    382 => "000000000000000000",
    383 => "000000000000000000",
    384 => "000000000000000000",
    385 => "000000000000000000",
    386 => "000000000000000000",
    387 => "000000000000000000",
    388 => "000000000000000000",
    389 => "000000000000000000",
    390 => "000000000000000000",
    391 => "000000000000000000",
    392 => "000000000000000000",
    393 => "000000000000000000",
    394 => "000000000000000000",
    395 => "000000000000000000",
    396 => "000000000000000000",
    397 => "000000000000000000",
    398 => "000000000000000000",
    399 => "000000000000000000",
    400 => "000000000000000000",
    401 => "000000000000000000",
    402 => "000000000000000000",
    403 => "000000000000000000",
    404 => "000000000000000000",
    405 => "000000000000000000",
    406 => "000000000000000000",
    407 => "000000000000000000",
    408 => "000000000000000000",
    409 => "000000000000000000",
    410 => "000000000000000000",
    411 => "000000000000000000",
    412 => "000000000000000000",
    413 => "000000000000000000",
    414 => "000000000000000000",
    415 => "000000000000000000",
    416 => "000000000000000000",
    417 => "000000000000000000",
    418 => "000000000000000000",
    419 => "000000000000000000",
    420 => "000000000000000000",
    421 => "000000000000000000",
    422 => "000000000000000000",
    423 => "000000000000000000",
    424 => "000000000000000000",
    425 => "000000000000000000",
    426 => "000000000000000000",
    427 => "000000000000000000",
    428 => "000000000000000000",
    429 => "000000000000000000",
    430 => "000000000000000000",
    431 => "000000000000000000",
    432 => "000000000000000000",
    433 => "000000000000000000",
    434 => "000000000000000000",
    435 => "000000000000000000",
    436 => "000000000000000000",
    437 => "000000000000000000",
    438 => "000000000000000000",
    439 => "000000000000000000",
    440 => "000000000000000000",
    441 => "000000000000000000",
    442 => "000000000000000000",
    443 => "000000000000000000",
    444 => "000000000000000000",
    445 => "000000000000000000",
    446 => "000000000000000000",
    447 => "000000000000000000",
    448 => "000000000000000000",
    449 => "000000000000000000",
    450 => "000000000000000000",
    451 => "000000000000000000",
    452 => "000000000000000000",
    453 => "000000000000000000",
    454 => "000000000000000000",
    455 => "000000000000000000",
    456 => "000000000000000000",
    457 => "000000000000000000",
    458 => "000000000000000000",
    459 => "000000000000000000",
    460 => "000000000000000000",
    461 => "000000000000000000",
    462 => "000000000000000000",
    463 => "000000000000000000",
    464 => "000000000000000000",
    465 => "000000000000000000",
    466 => "000000000000000000",
    467 => "000000000000000000",
    468 => "000000000000000000",
    469 => "000000000000000000",
    470 => "000000000000000000",
    471 => "000000000000000000",
    472 => "000000000000000000",
    473 => "000000000000000000",
    474 => "000000000000000000",
    475 => "000000000000000000",
    476 => "000000000000000000",
    477 => "000000000000000000",
    478 => "000000000000000000",
    479 => "000000000000000000",
    480 => "000000000000000000",
    481 => "000000000000000000",
    482 => "000000000000000000",
    483 => "000000000000000000",
    484 => "000000000000000000",
    485 => "000000000000000000",
    486 => "000000000000000000",
    487 => "000000000000000000",
    488 => "000000000000000000",
    489 => "000000000000000000",
    490 => "000000000000000000",
    491 => "000000000000000000",
    492 => "000000000000000000",
    493 => "000000000000000000",
    494 => "000000000000000000",
    495 => "000000000000000000",
    496 => "000000000000000000",
    497 => "000000000000000000",
    498 => "000000000000000000",
    499 => "000000000000000000",
    500 => "000000000000000000",
    501 => "000000000000000000",
    502 => "000000000000000000",
    503 => "000000000000000000",
    504 => "000000000000000000",
    505 => "000000000000000000",
    506 => "000000000000000000",
    507 => "000000000000000000",
    508 => "000000000000000000",
    509 => "000000000000000000",
    510 => "000000000000000000",
    511 => "000000000000000000",
    512 => "000000000000000000",
    513 => "000000000000000000",
    514 => "000000000000000000",
    515 => "000000000000000000",
    516 => "000000000000000000",
    517 => "000000000000000000",
    518 => "000000000000000000",
    519 => "000000000000000000",
    520 => "000000000000000000",
    521 => "000000000000000000",
    522 => "000000000000000000",
    523 => "000000000000000000",
    524 => "000000000000000000",
    525 => "000000000000000000",
    526 => "000000000000000000",
    527 => "000000000000000000",
    528 => "000000000000000000",
    529 => "000000000000000000",
    530 => "000000000000000000",
    531 => "000000000000000000",
    532 => "000000000000000000",
    533 => "000000000000000000",
    534 => "000000000000000000",
    535 => "000000000000000000",
    536 => "000000000000000000",
    537 => "000000000000000000",
    538 => "000000000000000000",
    539 => "000000000000000000",
    540 => "000000000000000000",
    541 => "000000000000000000",
    542 => "000000000000000000",
    543 => "000000000000000000",
    544 => "000000000000000000",
    545 => "000000000000000000",
    546 => "000000000000000000",
    547 => "000000000000000000",
    548 => "000000000000000000",
    549 => "000000000000000000",
    550 => "000000000000000000",
    551 => "000000000000000000",
    552 => "000000000000000000",
    553 => "000000000000000000",
    554 => "000000000000000000",
    555 => "000000000000000000",
    556 => "000000000000000000",
    557 => "000000000000000000",
    558 => "000000000000000000",
    559 => "000000000000000000",
    560 => "000000000000000000",
    561 => "000000000000000000",
    562 => "000000000000000000",
    563 => "000000000000000000",
    564 => "000000000000000000",
    565 => "000000000000000000",
    566 => "000000000000000000",
    567 => "000000000000000000",
    568 => "000000000000000000",
    569 => "000000000000000000",
    570 => "000000000000000000",
    571 => "000000000000000000",
    572 => "000000000000000000",
    573 => "000000000000000000",
    574 => "000000000000000000",
    575 => "000000000000000000",
    576 => "000000000000000000",
    577 => "000000000000000000",
    578 => "000000000000000000",
    579 => "000000000000000000",
    580 => "000000000000000000",
    581 => "000000000000000000",
    582 => "000000000000000000",
    583 => "000000000000000000",
    584 => "000000000000000000",
    585 => "000000000000000000",
    586 => "000000000000000000",
    587 => "000000000000000000",
    588 => "000000000000000000",
    589 => "000000000000000000",
    590 => "000000000000000000",
    591 => "000000000000000000",
    592 => "000000000000000000",
    593 => "000000000000000000",
    594 => "000000000000000000",
    595 => "000000000000000000",
    596 => "000000000000000000",
    597 => "000000000000000000",
    598 => "000000000000000000",
    599 => "000000000000000000",
    600 => "000000000000000000",
    601 => "000000000000000000",
    602 => "000000000000000000",
    603 => "000000000000000000",
    604 => "000000000000000000",
    605 => "000000000000000000",
    606 => "000000000000000000",
    607 => "000000000000000000",
    608 => "000000000000000000",
    609 => "000000000000000000",
    610 => "000000000000000000",
    611 => "000000000000000000",
    612 => "000000000000000000",
    613 => "000000000000000000",
    614 => "000000000000000000",
    615 => "000000000000000000",
    616 => "000000000000000000",
    617 => "000000000000000000",
    618 => "000000000000000000",
    619 => "000000000000000000",
    620 => "000000000000000000",
    621 => "000000000000000000",
    622 => "000000000000000000",
    623 => "000000000000000000",
    624 => "000000000000000000",
    625 => "000000000000000000",
    626 => "000000000000000000",
    627 => "000000000000000000",
    628 => "000000000000000000",
    629 => "000000000000000000",
    630 => "000000000000000000",
    631 => "000000000000000000",
    632 => "000000000000000000",
    633 => "000000000000000000",
    634 => "000000000000000000",
    635 => "000000000000000000",
    636 => "000000000000000000",
    637 => "000000000000000000",
    638 => "000000000000000000",
    639 => "000000000000000000",
    640 => "000000000000000000",
    641 => "000000000000000000",
    642 => "000000000000000000",
    643 => "000000000000000000",
    644 => "000000000000000000",
    645 => "000000000000000000",
    646 => "000000000000000000",
    647 => "000000000000000000",
    648 => "000000000000000000",
    649 => "000000000000000000",
    650 => "000000000000000000",
    651 => "000000000000000000",
    652 => "000000000000000000",
    653 => "000000000000000000",
    654 => "000000000000000000",
    655 => "000000000000000000",
    656 => "000000000000000000",
    657 => "000000000000000000",
    658 => "000000000000000000",
    659 => "000000000000000000",
    660 => "000000000000000000",
    661 => "000000000000000000",
    662 => "000000000000000000",
    663 => "000000000000000000",
    664 => "000000000000000000",
    665 => "000000000000000000",
    666 => "000000000000000000",
    667 => "000000000000000000",
    668 => "000000000000000000",
    669 => "000000000000000000",
    670 => "000000000000000000",
    671 => "000000000000000000",
    672 => "000000000000000000",
    673 => "000000000000000000",
    674 => "000000000000000000",
    675 => "000000000000000000",
    676 => "000000000000000000",
    677 => "000000000000000000",
    678 => "000000000000000000",
    679 => "000000000000000000",
    680 => "000000000000000000",
    681 => "000000000000000000",
    682 => "000000000000000000",
    683 => "000000000000000000",
    684 => "000000000000000000",
    685 => "000000000000000000",
    686 => "000000000000000000",
    687 => "000000000000000000",
    688 => "000000000000000000",
    689 => "000000000000000000",
    690 => "000000000000000000",
    691 => "000000000000000000",
    692 => "000000000000000000",
    693 => "000000000000000000",
    694 => "000000000000000000",
    695 => "000000000000000000",
    696 => "000000000000000000",
    697 => "000000000000000000",
    698 => "000000000000000000",
    699 => "000000000000000000",
    700 => "000000000000000000",
    701 => "000000000000000000",
    702 => "000000000000000000",
    703 => "000000000000000000",
    704 => "000000000000000000",
    705 => "000000000000000000",
    706 => "000000000000000000",
    707 => "000000000000000000",
    708 => "000000000000000000",
    709 => "000000000000000000",
    710 => "000000000000000000",
    711 => "000000000000000000",
    712 => "000000000000000000",
    713 => "000000000000000000",
    714 => "000000000000000000",
    715 => "000000000000000000",
    716 => "000000000000000000",
    717 => "000000000000000000",
    718 => "000000000000000000",
    719 => "000000000000000000",
    720 => "000000000000000000",
    721 => "000000000000000000",
    722 => "000000000000000000",
    723 => "000000000000000000",
    724 => "000000000000000000",
    725 => "000000000000000000",
    726 => "000000000000000000",
    727 => "000000000000000000",
    728 => "000000000000000000",
    729 => "000000000000000000",
    730 => "000000000000000000",
    731 => "000000000000000000",
    732 => "000000000000000000",
    733 => "000000000000000000",
    734 => "000000000000000000",
    735 => "000000000000000000",
    736 => "000000000000000000",
    737 => "000000000000000000",
    738 => "000000000000000000",
    739 => "000000000000000000",
    740 => "000000000000000000",
    741 => "000000000000000000",
    742 => "000000000000000000",
    743 => "000000000000000000",
    744 => "000000000000000000",
    745 => "000000000000000000",
    746 => "000000000000000000",
    747 => "000000000000000000",
    748 => "000000000000000000",
    749 => "000000000000000000",
    750 => "000000000000000000",
    751 => "000000000000000000",
    752 => "000000000000000000",
    753 => "000000000000000000",
    754 => "000000000000000000",
    755 => "000000000000000000",
    756 => "000000000000000000",
    757 => "000000000000000000",
    758 => "000000000000000000",
    759 => "000000000000000000",
    760 => "000000000000000000",
    761 => "000000000000000000",
    762 => "000000000000000000",
    763 => "000000000000000000",
    764 => "000000000000000000",
    765 => "000000000000000000",
    766 => "000000000000000000",
    767 => "000000000000000000",
    768 => "000000000000000000",
    769 => "000000000000000000",
    770 => "000000000000000000",
    771 => "000000000000000000",
    772 => "000000000000000000",
    773 => "000000000000000000",
    774 => "000000000000000000",
    775 => "000000000000000000",
    776 => "000000000000000000",
    777 => "000000000000000000",
    778 => "000000000000000000",
    779 => "000000000000000000",
    780 => "000000000000000000",
    781 => "000000000000000000",
    782 => "000000000000000000",
    783 => "000000000000000000",
    784 => "000000000000000000",
    785 => "000000000000000000",
    786 => "000000000000000000",
    787 => "000000000000000000",
    788 => "000000000000000000",
    789 => "000000000000000000",
    790 => "000000000000000000",
    791 => "000000000000000000",
    792 => "000000000000000000",
    793 => "000000000000000000",
    794 => "000000000000000000",
    795 => "000000000000000000",
    796 => "000000000000000000",
    797 => "000000000000000000",
    798 => "000000000000000000",
    799 => "000000000000000000",
    800 => "000000000000000000",
    801 => "000000000000000000",
    802 => "000000000000000000",
    803 => "000000000000000000",
    804 => "000000000000000000",
    805 => "000000000000000000",
    806 => "000000000000000000",
    807 => "000000000000000000",
    808 => "000000000000000000",
    809 => "000000000000000000",
    810 => "000000000000000000",
    811 => "000000000000000000",
    812 => "000000000000000000",
    813 => "000000000000000000",
    814 => "000000000000000000",
    815 => "000000000000000000",
    816 => "000000000000000000",
    817 => "000000000000000000",
    818 => "000000000000000000",
    819 => "000000000000000000",
    820 => "000000000000000000",
    821 => "000000000000000000",
    822 => "000000000000000000",
    823 => "000000000000000000",
    824 => "000000000000000000",
    825 => "000000000000000000",
    826 => "000000000000000000",
    827 => "000000000000000000",
    828 => "000000000000000000",
    829 => "000000000000000000",
    830 => "000000000000000000",
    831 => "000000000000000000",
    832 => "000000000000000000",
    833 => "000000000000000000",
    834 => "000000000000000000",
    835 => "000000000000000000",
    836 => "000000000000000000",
    837 => "000000000000000000",
    838 => "000000000000000000",
    839 => "000000000000000000",
    840 => "000000000000000000",
    841 => "000000000000000000",
    842 => "000000000000000000",
    843 => "000000000000000000",
    844 => "000000000000000000",
    845 => "000000000000000000",
    846 => "000000000000000000",
    847 => "000000000000000000",
    848 => "000000000000000000",
    849 => "000000000000000000",
    850 => "000000000000000000",
    851 => "000000000000000000",
    852 => "000000000000000000",
    853 => "000000000000000000",
    854 => "000000000000000000",
    855 => "000000000000000000",
    856 => "000000000000000000",
    857 => "000000000000000000",
    858 => "000000000000000000",
    859 => "000000000000000000",
    860 => "000000000000000000",
    861 => "000000000000000000",
    862 => "000000000000000000",
    863 => "000000000000000000",
    864 => "000000000000000000",
    865 => "000000000000000000",
    866 => "000000000000000000",
    867 => "000000000000000000",
    868 => "000000000000000000",
    869 => "000000000000000000",
    870 => "000000000000000000",
    871 => "000000000000000000",
    872 => "000000000000000000",
    873 => "000000000000000000",
    874 => "000000000000000000",
    875 => "000000000000000000",
    876 => "000000000000000000",
    877 => "000000000000000000",
    878 => "000000000000000000",
    879 => "000000000000000000",
    880 => "000000000000000000",
    881 => "000000000000000000",
    882 => "000000000000000000",
    883 => "000000000000000000",
    884 => "000000000000000000",
    885 => "000000000000000000",
    886 => "000000000000000000",
    887 => "000000000000000000",
    888 => "000000000000000000",
    889 => "000000000000000000",
    890 => "000000000000000000",
    891 => "000000000000000000",
    892 => "000000000000000000",
    893 => "000000000000000000",
    894 => "000000000000000000",
    895 => "000000000000000000",
    896 => "000000000000000000",
    897 => "000000000000000000",
    898 => "000000000000000000",
    899 => "000000000000000000",
    900 => "000000000000000000",
    901 => "000000000000000000",
    902 => "000000000000000000",
    903 => "000000000000000000",
    904 => "000000000000000000",
    905 => "000000000000000000",
    906 => "000000000000000000",
    907 => "000000000000000000",
    908 => "000000000000000000",
    909 => "000000000000000000",
    910 => "000000000000000000",
    911 => "000000000000000000",
    912 => "000000000000000000",
    913 => "000000000000000000",
    914 => "000000000000000000",
    915 => "000000000000000000",
    916 => "000000000000000000",
    917 => "000000000000000000",
    918 => "000000000000000000",
    919 => "000000000000000000",
    920 => "000000000000000000",
    921 => "000000000000000000",
    922 => "000000000000000000",
    923 => "000000000000000000",
    924 => "000000000000000000",
    925 => "000000000000000000",
    926 => "000000000000000000",
    927 => "000000000000000000",
    928 => "000000000000000000",
    929 => "000000000000000000",
    930 => "000000000000000000",
    931 => "000000000000000000",
    932 => "000000000000000000",
    933 => "000000000000000000",
    934 => "000000000000000000",
    935 => "000000000000000000",
    936 => "000000000000000000",
    937 => "000000000000000000",
    938 => "000000000000000000",
    939 => "000000000000000000",
    940 => "000000000000000000",
    941 => "000000000000000000",
    942 => "000000000000000000",
    943 => "000000000000000000",
    944 => "000000000000000000",
    945 => "000000000000000000",
    946 => "000000000000000000",
    947 => "000000000000000000",
    948 => "000000000000000000",
    949 => "000000000000000000",
    950 => "000000000000000000",
    951 => "000000000000000000",
    952 => "000000000000000000",
    953 => "000000000000000000",
    954 => "000000000000000000",
    955 => "000000000000000000",
    956 => "000000000000000000",
    957 => "000000000000000000",
    958 => "000000000000000000",
    959 => "000000000000000000",
    960 => "000000000000000000",
    961 => "000000000000000000",
    962 => "000000000000000000",
    963 => "000000000000000000",
    964 => "000000000000000000",
    965 => "000000000000000000",
    966 => "000000000000000000",
    967 => "000000000000000000",
    968 => "000000000000000000",
    969 => "000000000000000000",
    970 => "000000000000000000",
    971 => "000000000000000000",
    972 => "000000000000000000",
    973 => "000000000000000000",
    974 => "000000000000000000",
    975 => "000000000000000000",
    976 => "000000000000000000",
    977 => "000000000000000000",
    978 => "000000000000000000",
    979 => "000000000000000000",
    980 => "000000000000000000",
    981 => "000000000000000000",
    982 => "000000000000000000",
    983 => "000000000000000000",
    984 => "000000000000000000",
    985 => "000000000000000000",
    986 => "000000000000000000",
    987 => "000000000000000000",
    988 => "000000000000000000",
    989 => "000000000000000000",
    990 => "000000000000000000",
    991 => "000000000000000000",
    992 => "000000000000000000",
    993 => "000000000000000000",
    994 => "000000000000000000",
    995 => "000000000000000000",
    996 => "000000000000000000",
    997 => "000000000000000000",
    998 => "000000000000000000",
    999 => "000000000000000000",
    1000 => "000000000000000000",
    1001 => "000000000000000000",
    1002 => "000000000000000000",
    1003 => "000000000000000000",
    1004 => "000000000000000000",
    1005 => "000000000000000000",
    1006 => "000000000000000000",
    1007 => "000000000000000000",
    1008 => "000000000000000000",
    1009 => "000000000000000000",
    1010 => "000000000000000000",
    1011 => "000000000000000000",
    1012 => "000000000000000000",
    1013 => "000000000000000000",
    1014 => "000000000000000000",
    1015 => "000000000000000000",
    1016 => "000000000000000000",
    1017 => "000000000000000000",
    1018 => "000000000000000000",
    1019 => "000000000000000000",
    1020 => "000000000000000000",
    1021 => "000000000000000000",
    1022 => "000000000000000000",
    1023 => "000000000000000000",
    1024 => "000000000000000000",
    1025 => "000000000000000000",
    1026 => "000000000000000000",
    1027 => "000000000000000000",
    1028 => "000000000000000000",
    1029 => "000000000000000000",
    1030 => "000000000000000000",
    1031 => "000000000000000000",
    1032 => "000000000000000000",
    1033 => "000000000000000000",
    1034 => "000000000000000000",
    1035 => "000000000000000000",
    1036 => "000000000000000000",
    1037 => "000000000000000000",
    1038 => "000000000000000000",
    1039 => "000000000000000000",
    1040 => "000000000000000000",
    1041 => "000000000000000000",
    1042 => "000000000000000000",
    1043 => "000000000000000000",
    1044 => "000000000000000000",
    1045 => "000000000000000000",
    1046 => "000000000000000000",
    1047 => "000000000000000000",
    1048 => "000000000000000000",
    1049 => "000000000000000000",
    1050 => "000000000000000000",
    1051 => "000000000000000000",
    1052 => "000000000000000000",
    1053 => "000000000000000000",
    1054 => "000000000000000000",
    1055 => "000000000000000000",
    1056 => "000000000000000000",
    1057 => "000000000000000000",
    1058 => "000000000000000000",
    1059 => "000000000000000000",
    1060 => "000000000000000000",
    1061 => "000000000000000000",
    1062 => "000000000000000000",
    1063 => "000000000000000000",
    1064 => "000000000000000000",
    1065 => "000000000000000000",
    1066 => "000000000000000000",
    1067 => "000000000000000000",
    1068 => "000000000000000000",
    1069 => "000000000000000000",
    1070 => "000000000000000000",
    1071 => "000000000000000000",
    1072 => "000000000000000000",
    1073 => "000000000000000000",
    1074 => "000000000000000000",
    1075 => "000000000000000000",
    1076 => "000000000000000000",
    1077 => "000000000000000000",
    1078 => "000000000000000000",
    1079 => "000000000000000000",
    1080 => "000000000000000000",
    1081 => "000000000000000000",
    1082 => "000000000000000000",
    1083 => "000000000000000000",
    1084 => "000000000000000000",
    1085 => "000000000000000000",
    1086 => "000000000000000000",
    1087 => "000000000000000000",
    1088 => "000000000000000000",
    1089 => "000000000000000000",
    1090 => "000000000000000000",
    1091 => "000000000000000000",
    1092 => "000000000000000000",
    1093 => "000000000000000000",
    1094 => "000000000000000000",
    1095 => "000000000000000000",
    1096 => "000000000000000000",
    1097 => "000000000000000000",
    1098 => "000000000000000000",
    1099 => "000000000000000000",
    1100 => "000000000000000000",
    1101 => "000000000000000000",
    1102 => "000000000000000000",
    1103 => "000000000000000000",
    1104 => "000000000000000000",
    1105 => "000000000000000000",
    1106 => "000000000000000000",
    1107 => "000000000000000000",
    1108 => "000000000000000000",
    1109 => "000000000000000000",
    1110 => "000000000000000000",
    1111 => "000000000000000000",
    1112 => "000000000000000000",
    1113 => "000000000000000000",
    1114 => "000000000000000000",
    1115 => "000000000000000000",
    1116 => "000000000000000000",
    1117 => "000000000000000000",
    1118 => "000000000000000000",
    1119 => "000000000000000000",
    1120 => "000000000000000000",
    1121 => "000000000000000000",
    1122 => "000000000000000000",
    1123 => "000000000000000000",
    1124 => "000000000000000000",
    1125 => "000000000000000000",
    1126 => "000000000000000000",
    1127 => "000000000000000000",
    1128 => "000000000000000000",
    1129 => "000000000000000000",
    1130 => "000000000000000000",
    1131 => "000000000000000000",
    1132 => "000000000000000000",
    1133 => "000000000000000000",
    1134 => "000000000000000000",
    1135 => "000000000000000000",
    1136 => "000000000000000000",
    1137 => "000000000000000000",
    1138 => "000000000000000000",
    1139 => "000000000000000000",
    1140 => "000000000000000000",
    1141 => "000000000000000000",
    1142 => "000000000000000000",
    1143 => "000000000000000000",
    1144 => "000000000000000000",
    1145 => "000000000000000000",
    1146 => "000000000000000000",
    1147 => "000000000000000000",
    1148 => "000000000000000000",
    1149 => "000000000000000000",
    1150 => "000000000000000000",
    1151 => "000000000000000000",
    1152 => "000000000000000000",
    1153 => "000000000000000000",
    1154 => "000000000000000000",
    1155 => "000000000000000000",
    1156 => "000000000000000000",
    1157 => "000000000000000000",
    1158 => "000000000000000000",
    1159 => "000000000000000000",
    1160 => "000000000000000000",
    1161 => "000000000000000000",
    1162 => "000000000000000000",
    1163 => "000000000000000000",
    1164 => "000000000000000000",
    1165 => "000000000000000000",
    1166 => "000000000000000000",
    1167 => "000000000000000000",
    1168 => "000000000000000000",
    1169 => "000000000000000000",
    1170 => "000000000000000000",
    1171 => "000000000000000000",
    1172 => "000000000000000000",
    1173 => "000000000000000000",
    1174 => "000000000000000000",
    1175 => "000000000000000000",
    1176 => "000000000000000000",
    1177 => "000000000000000000",
    1178 => "000000000000000000",
    1179 => "000000000000000000",
    1180 => "000000000000000000",
    1181 => "000000000000000000",
    1182 => "000000000000000000",
    1183 => "000000000000000000",
    1184 => "000000000000000000",
    1185 => "000000000000000000",
    1186 => "000000000000000000",
    1187 => "000000000000000000",
    1188 => "000000000000000000",
    1189 => "000000000000000000",
    1190 => "000000000000000000",
    1191 => "000000000000000000",
    1192 => "000000000000000000",
    1193 => "000000000000000000",
    1194 => "000000000000000000",
    1195 => "000000000000000000",
    1196 => "000000000000000000",
    1197 => "000000000000000000",
    1198 => "000000000000000000",
    1199 => "000000000000000000",
    1200 => "000000000000000000",
    1201 => "000000000000000000",
    1202 => "000000000000000000",
    1203 => "000000000000000000",
    1204 => "000000000000000000",
    1205 => "000000000000000000",
    1206 => "000000000000000000",
    1207 => "000000000000000000",
    1208 => "000000000000000000",
    1209 => "000000000000000000",
    1210 => "000000000000000000",
    1211 => "000000000000000000",
    1212 => "000000000000000000",
    1213 => "000000000000000000",
    1214 => "000000000000000000",
    1215 => "000000000000000000",
    1216 => "000000000000000000",
    1217 => "000000000000000000",
    1218 => "000000000000000000",
    1219 => "000000000000000000",
    1220 => "000000000000000000",
    1221 => "000000000000000000",
    1222 => "000000000000000000",
    1223 => "000000000000000000",
    1224 => "000000000000000000",
    1225 => "000000000000000000",
    1226 => "000000000000000000",
    1227 => "000000000000000000",
    1228 => "000000000000000000",
    1229 => "000000000000000000",
    1230 => "000000000000000000",
    1231 => "000000000000000000",
    1232 => "000000000000000000",
    1233 => "000000000000000000",
    1234 => "000000000000000000",
    1235 => "000000000000000000",
    1236 => "000000000000000000",
    1237 => "000000000000000000",
    1238 => "000000000000000000",
    1239 => "000000000000000000",
    1240 => "000000000000000000",
    1241 => "000000000000000000",
    1242 => "000000000000000000",
    1243 => "000000000000000000",
    1244 => "000000000000000000",
    1245 => "000000000000000000",
    1246 => "000000000000000000",
    1247 => "000000000000000000",
    1248 => "000000000000000000",
    1249 => "000000000000000000",
    1250 => "000000000000000000",
    1251 => "000000000000000000",
    1252 => "000000000000000000",
    1253 => "000000000000000000",
    1254 => "000000000000000000",
    1255 => "000000000000000000",
    1256 => "000000000000000000",
    1257 => "000000000000000000",
    1258 => "000000000000000000",
    1259 => "000000000000000000",
    1260 => "000000000000000000",
    1261 => "000000000000000000",
    1262 => "000000000000000000",
    1263 => "000000000000000000",
    1264 => "000000000000000000",
    1265 => "000000000000000000",
    1266 => "000000000000000000",
    1267 => "000000000000000000",
    1268 => "000000000000000000",
    1269 => "000000000000000000",
    1270 => "000000000000000000",
    1271 => "000000000000000000",
    1272 => "000000000000000000",
    1273 => "000000000000000000",
    1274 => "000000000000000000",
    1275 => "000000000000000000",
    1276 => "000000000000000000",
    1277 => "000000000000000000",
    1278 => "000000000000000000",
    1279 => "000000000000000000",
    1280 => "000000000000000000",
    1281 => "000000000000000000",
    1282 => "000000000000000000",
    1283 => "000000000000000000",
    1284 => "000000000000000000",
    1285 => "000000000000000000",
    1286 => "000000000000000000",
    1287 => "000000000000000000",
    1288 => "000000000000000000",
    1289 => "000000000000000000",
    1290 => "000000000000000000",
    1291 => "000000000000000000",
    1292 => "000000000000000000",
    1293 => "000000000000000000",
    1294 => "000000000000000000",
    1295 => "000000000000000000",
    1296 => "000000000000000000",
    1297 => "000000000000000000",
    1298 => "000000000000000000",
    1299 => "000000000000000000",
    1300 => "000000000000000000",
    1301 => "000000000000000000",
    1302 => "000000000000000000",
    1303 => "000000000000000000",
    1304 => "000000000000000000",
    1305 => "000000000000000000",
    1306 => "000000000000000000",
    1307 => "000000000000000000",
    1308 => "000000000000000000",
    1309 => "000000000000000000",
    1310 => "000000000000000000",
    1311 => "000000000000000000",
    1312 => "000000000000000000",
    1313 => "000000000000000000",
    1314 => "000000000000000000",
    1315 => "000000000000000000",
    1316 => "000000000000000000",
    1317 => "000000000000000000",
    1318 => "000000000000000000",
    1319 => "000000000000000000",
    1320 => "000000000000000000",
    1321 => "000000000000000000",
    1322 => "000000000000000000",
    1323 => "000000000000000000",
    1324 => "000000000000000000",
    1325 => "000000000000000000",
    1326 => "000000000000000000",
    1327 => "000000000000000000",
    1328 => "000000000000000000",
    1329 => "000000000000000000",
    1330 => "000000000000000000",
    1331 => "000000000000000000",
    1332 => "000000000000000000",
    1333 => "000000000000000000",
    1334 => "000000000000000000",
    1335 => "000000000000000000",
    1336 => "000000000000000000",
    1337 => "000000000000000000",
    1338 => "000000000000000000",
    1339 => "000000000000000000",
    1340 => "000000000000000000",
    1341 => "000000000000000000",
    1342 => "000000000000000000",
    1343 => "000000000000000000",
    1344 => "000000000000000000",
    1345 => "000000000000000000",
    1346 => "000000000000000000",
    1347 => "000000000000000000",
    1348 => "000000000000000000",
    1349 => "000000000000000000",
    1350 => "000000000000000000",
    1351 => "000000000000000000",
    1352 => "000000000000000000",
    1353 => "000000000000000000",
    1354 => "000000000000000000",
    1355 => "000000000000000000",
    1356 => "000000000000000000",
    1357 => "000000000000000000",
    1358 => "000000000000000000",
    1359 => "000000000000000000",
    1360 => "000000000000000000",
    1361 => "000000000000000000",
    1362 => "000000000000000000",
    1363 => "000000000000000000",
    1364 => "000000000000000000",
    1365 => "000000000000000000",
    1366 => "000000000000000000",
    1367 => "000000000000000000",
    1368 => "000000000000000000",
    1369 => "000000000000000000",
    1370 => "000000000000000000",
    1371 => "000000000000000000",
    1372 => "000000000000000000",
    1373 => "000000000000000000",
    1374 => "000000000000000000",
    1375 => "000000000000000000",
    1376 => "000000000000000000",
    1377 => "000000000000000000",
    1378 => "000000000000000000",
    1379 => "000000000000000000",
    1380 => "000000000000000000",
    1381 => "000000000000000000",
    1382 => "000000000000000000",
    1383 => "000000000000000000",
    1384 => "000000000000000000",
    1385 => "000000000000000000",
    1386 => "000000000000000000",
    1387 => "000000000000000000",
    1388 => "000000000000000000",
    1389 => "000000000000000000",
    1390 => "000000000000000000",
    1391 => "000000000000000000",
    1392 => "000000000000000000",
    1393 => "000000000000000000",
    1394 => "000000000000000000",
    1395 => "000000000000000000",
    1396 => "000000000000000000",
    1397 => "000000000000000000",
    1398 => "000000000000000000",
    1399 => "000000000000000000",
    1400 => "000000000000000000",
    1401 => "000000000000000000",
    1402 => "000000000000000000",
    1403 => "000000000000000000",
    1404 => "000000000000000000",
    1405 => "000000000000000000",
    1406 => "000000000000000000",
    1407 => "000000000000000000",
    1408 => "000000000000000000",
    1409 => "000000000000000000",
    1410 => "000000000000000000",
    1411 => "000000000000000000",
    1412 => "000000000000000000",
    1413 => "000000000000000000",
    1414 => "000000000000000000",
    1415 => "000000000000000000",
    1416 => "000000000000000000",
    1417 => "000000000000000000",
    1418 => "000000000000000000",
    1419 => "000000000000000000",
    1420 => "000000000000000000",
    1421 => "000000000000000000",
    1422 => "000000000000000000",
    1423 => "000000000000000000",
    1424 => "000000000000000000",
    1425 => "000000000000000000",
    1426 => "000000000000000000",
    1427 => "000000000000000000",
    1428 => "000000000000000000",
    1429 => "000000000000000000",
    1430 => "000000000000000000",
    1431 => "000000000000000000",
    1432 => "000000000000000000",
    1433 => "000000000000000000",
    1434 => "000000000000000000",
    1435 => "000000000000000000",
    1436 => "000000000000000000",
    1437 => "000000000000000000",
    1438 => "000000000000000000",
    1439 => "000000000000000000",
    1440 => "000000000000000000",
    1441 => "000000000000000000",
    1442 => "000000000000000000",
    1443 => "000000000000000000",
    1444 => "000000000000000000",
    1445 => "000000000000000000",
    1446 => "000000000000000000",
    1447 => "000000000000000000",
    1448 => "000000000000000000",
    1449 => "000000000000000000",
    1450 => "000000000000000000",
    1451 => "000000000000000000",
    1452 => "000000000000000000",
    1453 => "000000000000000000",
    1454 => "000000000000000000",
    1455 => "000000000000000000",
    1456 => "000000000000000000",
    1457 => "000000000000000000",
    1458 => "000000000000000000",
    1459 => "000000000000000000",
    1460 => "000000000000000000",
    1461 => "000000000000000000",
    1462 => "000000000000000000",
    1463 => "000000000000000000",
    1464 => "000000000000000000",
    1465 => "000000000000000000",
    1466 => "000000000000000000",
    1467 => "000000000000000000",
    1468 => "000000000000000000",
    1469 => "000000000000000000",
    1470 => "000000000000000000",
    1471 => "000000000000000000",
    1472 => "000000000000000000",
    1473 => "000000000000000000",
    1474 => "000000000000000000",
    1475 => "000000000000000000",
    1476 => "000000000000000000",
    1477 => "000000000000000000",
    1478 => "000000000000000000",
    1479 => "000000000000000000",
    1480 => "000000000000000000",
    1481 => "000000000000000000",
    1482 => "000000000000000000",
    1483 => "000000000000000000",
    1484 => "000000000000000000",
    1485 => "000000000000000000",
    1486 => "000000000000000000",
    1487 => "000000000000000000",
    1488 => "000000000000000000",
    1489 => "000000000000000000",
    1490 => "000000000000000000",
    1491 => "000000000000000000",
    1492 => "000000000000000000",
    1493 => "000000000000000000",
    1494 => "000000000000000000",
    1495 => "000000000000000000",
    1496 => "000000000000000000",
    1497 => "000000000000000000",
    1498 => "000000000000000000",
    1499 => "000000000000000000",
    1500 => "000000000000000000",
    1501 => "000000000000000000",
    1502 => "000000000000000000",
    1503 => "000000000000000000",
    1504 => "000000000000000000",
    1505 => "000000000000000000",
    1506 => "000000000000000000",
    1507 => "000000000000000000",
    1508 => "000000000000000000",
    1509 => "000000000000000000",
    1510 => "000000000000000000",
    1511 => "000000000000000000",
    1512 => "000000000000000000",
    1513 => "000000000000000000",
    1514 => "000000000000000000",
    1515 => "000000000000000000",
    1516 => "000000000000000000",
    1517 => "000000000000000000",
    1518 => "000000000000000000",
    1519 => "000000000000000000",
    1520 => "000000000000000000",
    1521 => "000000000000000000",
    1522 => "000000000000000000",
    1523 => "000000000000000000",
    1524 => "000000000000000000",
    1525 => "000000000000000000",
    1526 => "000000000000000000",
    1527 => "000000000000000000",
    1528 => "000000000000000000",
    1529 => "000000000000000000",
    1530 => "000000000000000000",
    1531 => "000000000000000000",
    1532 => "000000000000000000",
    1533 => "000000000000000000",
    1534 => "000000000000000000",
    1535 => "000000000000000000",
    1536 => "000000000000000000",
    1537 => "000000000000000000",
    1538 => "000000000000000000",
    1539 => "000000000000000000",
    1540 => "000000000000000000",
    1541 => "000000000000000000",
    1542 => "000000000000000000",
    1543 => "000000000000000000",
    1544 => "000000000000000000",
    1545 => "000000000000000000",
    1546 => "000000000000000000",
    1547 => "000000000000000000",
    1548 => "000000000000000000",
    1549 => "000000000000000000",
    1550 => "000000000000000000",
    1551 => "000000000000000000",
    1552 => "000000000000000000",
    1553 => "000000000000000000",
    1554 => "000000000000000000",
    1555 => "000000000000000000",
    1556 => "000000000000000000",
    1557 => "000000000000000000",
    1558 => "000000000000000000",
    1559 => "000000000000000000",
    1560 => "000000000000000000",
    1561 => "000000000000000000",
    1562 => "000000000000000000",
    1563 => "000000000000000000",
    1564 => "000000000000000000",
    1565 => "000000000000000000",
    1566 => "000000000000000000",
    1567 => "000000000000000000",
    1568 => "000000000000000000",
    1569 => "000000000000000000",
    1570 => "000000000000000000",
    1571 => "000000000000000000",
    1572 => "000000000000000000",
    1573 => "000000000000000000",
    1574 => "000000000000000000",
    1575 => "000000000000000000",
    1576 => "000000000000000000",
    1577 => "000000000000000000",
    1578 => "000000000000000000",
    1579 => "000000000000000000",
    1580 => "000000000000000000",
    1581 => "000000000000000000",
    1582 => "000000000000000000",
    1583 => "000000000000000000",
    1584 => "000000000000000000",
    1585 => "000000000000000000",
    1586 => "000000000000000000",
    1587 => "000000000000000000",
    1588 => "000000000000000000",
    1589 => "000000000000000000",
    1590 => "000000000000000000",
    1591 => "000000000000000000",
    1592 => "000000000000000000",
    1593 => "000000000000000000",
    1594 => "000000000000000000",
    1595 => "000000000000000000",
    1596 => "000000000000000000",
    1597 => "000000000000000000",
    1598 => "000000000000000000",
    1599 => "000000000000000000",
    1600 => "000000000000000000",
    1601 => "000000000000000000",
    1602 => "000000000000000000",
    1603 => "000000000000000000",
    1604 => "000000000000000000",
    1605 => "000000000000000000",
    1606 => "000000000000000000",
    1607 => "000000000000000000",
    1608 => "000000000000000000",
    1609 => "000000000000000000",
    1610 => "000000000000000000",
    1611 => "000000000000000000",
    1612 => "000000000000000000",
    1613 => "000000000000000000",
    1614 => "000000000000000000",
    1615 => "000000000000000000",
    1616 => "000000000000000000",
    1617 => "000000000000000000",
    1618 => "000000000000000000",
    1619 => "000000000000000000",
    1620 => "000000000000000000",
    1621 => "000000000000000000",
    1622 => "000000000000000000",
    1623 => "000000000000000000",
    1624 => "000000000000000000",
    1625 => "000000000000000000",
    1626 => "000000000000000000",
    1627 => "000000000000000000",
    1628 => "000000000000000000",
    1629 => "000000000000000000",
    1630 => "000000000000000000",
    1631 => "000000000000000000",
    1632 => "000000000000000000",
    1633 => "000000000000000000",
    1634 => "000000000000000000",
    1635 => "000000000000000000",
    1636 => "000000000000000000",
    1637 => "000000000000000000",
    1638 => "000000000000000000",
    1639 => "000000000000000000",
    1640 => "000000000000000000",
    1641 => "000000000000000000",
    1642 => "000000000000000000",
    1643 => "000000000000000000",
    1644 => "000000000000000000",
    1645 => "000000000000000000",
    1646 => "000000000000000000",
    1647 => "000000000000000000",
    1648 => "000000000000000000",
    1649 => "000000000000000000",
    1650 => "000000000000000000",
    1651 => "000000000000000000",
    1652 => "000000000000000000",
    1653 => "000000000000000000",
    1654 => "000000000000000000",
    1655 => "000000000000000000",
    1656 => "000000000000000000",
    1657 => "000000000000000000",
    1658 => "000000000000000000",
    1659 => "000000000000000000",
    1660 => "000000000000000000",
    1661 => "000000000000000000",
    1662 => "000000000000000000",
    1663 => "000000000000000000",
    1664 => "000000000000000000",
    1665 => "000000000000000000",
    1666 => "000000000000000000",
    1667 => "000000000000000000",
    1668 => "000000000000000000",
    1669 => "000000000000000000",
    1670 => "000000000000000000",
    1671 => "000000000000000000",
    1672 => "000000000000000000",
    1673 => "000000000000000000",
    1674 => "000000000000000000",
    1675 => "000000000000000000",
    1676 => "000000000000000000",
    1677 => "000000000000000000",
    1678 => "000000000000000000",
    1679 => "000000000000000000",
    1680 => "000000000000000000",
    1681 => "000000000000000000",
    1682 => "000000000000000000",
    1683 => "000000000000000000",
    1684 => "000000000000000000",
    1685 => "000000000000000000",
    1686 => "000000000000000000",
    1687 => "000000000000000000",
    1688 => "000000000000000000",
    1689 => "000000000000000000",
    1690 => "000000000000000000",
    1691 => "000000000000000000",
    1692 => "000000000000000000",
    1693 => "000000000000000000",
    1694 => "000000000000000000",
    1695 => "000000000000000000",
    1696 => "000000000000000000",
    1697 => "000000000000000000",
    1698 => "000000000000000000",
    1699 => "000000000000000000",
    1700 => "000000000000000000",
    1701 => "000000000000000000",
    1702 => "000000000000000000",
    1703 => "000000000000000000",
    1704 => "000000000000000000",
    1705 => "000000000000000000",
    1706 => "000000000000000000",
    1707 => "000000000000000000",
    1708 => "000000000000000000",
    1709 => "000000000000000000",
    1710 => "000000000000000000",
    1711 => "000000000000000000",
    1712 => "000000000000000000",
    1713 => "000000000000000000",
    1714 => "000000000000000000",
    1715 => "000000000000000000",
    1716 => "000000000000000000",
    1717 => "000000000000000000",
    1718 => "000000000000000000",
    1719 => "000000000000000000",
    1720 => "000000000000000000",
    1721 => "000000000000000000",
    1722 => "000000000000000000",
    1723 => "000000000000000000",
    1724 => "000000000000000000",
    1725 => "000000000000000000",
    1726 => "000000000000000000",
    1727 => "000000000000000000",
    1728 => "000000000000000000",
    1729 => "000000000000000000",
    1730 => "000000000000000000",
    1731 => "000000000000000000",
    1732 => "000000000000000000",
    1733 => "000000000000000000",
    1734 => "000000000000000000",
    1735 => "000000000000000000",
    1736 => "000000000000000000",
    1737 => "000000000000000000",
    1738 => "000000000000000000",
    1739 => "000000000000000000",
    1740 => "000000000000000000",
    1741 => "000000000000000000",
    1742 => "000000000000000000",
    1743 => "000000000000000000",
    1744 => "000000000000000000",
    1745 => "000000000000000000",
    1746 => "000000000000000000",
    1747 => "000000000000000000",
    1748 => "000000000000000000",
    1749 => "000000000000000000",
    1750 => "000000000000000000",
    1751 => "000000000000000000",
    1752 => "000000000000000000",
    1753 => "000000000000000000",
    1754 => "000000000000000000",
    1755 => "000000000000000000",
    1756 => "000000000000000000",
    1757 => "000000000000000000",
    1758 => "000000000000000000",
    1759 => "000000000000000000",
    1760 => "000000000000000000",
    1761 => "000000000000000000",
    1762 => "000000000000000000",
    1763 => "000000000000000000",
    1764 => "000000000000000000",
    1765 => "000000000000000000",
    1766 => "000000000000000000",
    1767 => "000000000000000000",
    1768 => "000000000000000000",
    1769 => "000000000000000000",
    1770 => "000000000000000000",
    1771 => "000000000000000000",
    1772 => "000000000000000000",
    1773 => "000000000000000000",
    1774 => "000000000000000000",
    1775 => "000000000000000000",
    1776 => "000000000000000000",
    1777 => "000000000000000000",
    1778 => "000000000000000000",
    1779 => "000000000000000000",
    1780 => "000000000000000000",
    1781 => "000000000000000000",
    1782 => "000000000000000000",
    1783 => "000000000000000000",
    1784 => "000000000000000000",
    1785 => "000000000000000000",
    1786 => "000000000000000000",
    1787 => "000000000000000000",
    1788 => "000000000000000000",
    1789 => "000000000000000000",
    1790 => "000000000000000000",
    1791 => "000000000000000000",
    1792 => "000000000000000000",
    1793 => "000000000000000000",
    1794 => "000000000000000000",
    1795 => "000000000000000000",
    1796 => "000000000000000000",
    1797 => "000000000000000000",
    1798 => "000000000000000000",
    1799 => "000000000000000000",
    1800 => "000000000000000000",
    1801 => "000000000000000000",
    1802 => "000000000000000000",
    1803 => "000000000000000000",
    1804 => "000000000000000000",
    1805 => "000000000000000000",
    1806 => "000000000000000000",
    1807 => "000000000000000000",
    1808 => "000000000000000000",
    1809 => "000000000000000000",
    1810 => "000000000000000000",
    1811 => "000000000000000000",
    1812 => "000000000000000000",
    1813 => "000000000000000000",
    1814 => "000000000000000000",
    1815 => "000000000000000000",
    1816 => "000000000000000000",
    1817 => "000000000000000000",
    1818 => "000000000000000000",
    1819 => "000000000000000000",
    1820 => "000000000000000000",
    1821 => "000000000000000000",
    1822 => "000000000000000000",
    1823 => "000000000000000000",
    1824 => "000000000000000000",
    1825 => "000000000000000000",
    1826 => "000000000000000000",
    1827 => "000000000000000000",
    1828 => "000000000000000000",
    1829 => "000000000000000000",
    1830 => "000000000000000000",
    1831 => "000000000000000000",
    1832 => "000000000000000000",
    1833 => "000000000000000000",
    1834 => "000000000000000000",
    1835 => "000000000000000000",
    1836 => "000000000000000000",
    1837 => "000000000000000000",
    1838 => "000000000000000000",
    1839 => "000000000000000000",
    1840 => "000000000000000000",
    1841 => "000000000000000000",
    1842 => "000000000000000000",
    1843 => "000000000000000000",
    1844 => "000000000000000000",
    1845 => "000000000000000000",
    1846 => "000000000000000000",
    1847 => "000000000000000000",
    1848 => "000000000000000000",
    1849 => "000000000000000000",
    1850 => "000000000000000000",
    1851 => "000000000000000000",
    1852 => "000000000000000000",
    1853 => "000000000000000000",
    1854 => "000000000000000000",
    1855 => "000000000000000000",
    1856 => "000000000000000000",
    1857 => "000000000000000000",
    1858 => "000000000000000000",
    1859 => "000000000000000000",
    1860 => "000000000000000000",
    1861 => "000000000000000000",
    1862 => "000000000000000000",
    1863 => "000000000000000000",
    1864 => "000000000000000000",
    1865 => "000000000000000000",
    1866 => "000000000000000000",
    1867 => "000000000000000000",
    1868 => "000000000000000000",
    1869 => "000000000000000000",
    1870 => "000000000000000000",
    1871 => "000000000000000000",
    1872 => "000000000000000000",
    1873 => "000000000000000000",
    1874 => "000000000000000000",
    1875 => "000000000000000000",
    1876 => "000000000000000000",
    1877 => "000000000000000000",
    1878 => "000000000000000000",
    1879 => "000000000000000000",
    1880 => "000000000000000000",
    1881 => "000000000000000000",
    1882 => "000000000000000000",
    1883 => "000000000000000000",
    1884 => "000000000000000000",
    1885 => "000000000000000000",
    1886 => "000000000000000000",
    1887 => "000000000000000000",
    1888 => "000000000000000000",
    1889 => "000000000000000000",
    1890 => "000000000000000000",
    1891 => "000000000000000000",
    1892 => "000000000000000000",
    1893 => "000000000000000000",
    1894 => "000000000000000000",
    1895 => "000000000000000000",
    1896 => "000000000000000000",
    1897 => "000000000000000000",
    1898 => "000000000000000000",
    1899 => "000000000000000000",
    1900 => "000000000000000000",
    1901 => "000000000000000000",
    1902 => "000000000000000000",
    1903 => "000000000000000000",
    1904 => "000000000000000000",
    1905 => "000000000000000000",
    1906 => "000000000000000000",
    1907 => "000000000000000000",
    1908 => "000000000000000000",
    1909 => "000000000000000000",
    1910 => "000000000000000000",
    1911 => "000000000000000000",
    1912 => "000000000000000000",
    1913 => "000000000000000000",
    1914 => "000000000000000000",
    1915 => "000000000000000000",
    1916 => "000000000000000000",
    1917 => "000000000000000000",
    1918 => "000000000000000000",
    1919 => "000000000000000000",
    1920 => "000000000000000000",
    1921 => "000000000000000000",
    1922 => "000000000000000000",
    1923 => "000000000000000000",
    1924 => "000000000000000000",
    1925 => "000000000000000000",
    1926 => "000000000000000000",
    1927 => "000000000000000000",
    1928 => "000000000000000000",
    1929 => "000000000000000000",
    1930 => "000000000000000000",
    1931 => "000000000000000000",
    1932 => "000000000000000000",
    1933 => "000000000000000000",
    1934 => "000000000000000000",
    1935 => "000000000000000000",
    1936 => "000000000000000000",
    1937 => "000000000000000000",
    1938 => "000000000000000000",
    1939 => "000000000000000000",
    1940 => "000000000000000000",
    1941 => "000000000000000000",
    1942 => "000000000000000000",
    1943 => "000000000000000000",
    1944 => "000000000000000000",
    1945 => "000000000000000000",
    1946 => "000000000000000000",
    1947 => "000000000000000000",
    1948 => "000000000000000000",
    1949 => "000000000000000000",
    1950 => "000000000000000000",
    1951 => "000000000000000000",
    1952 => "000000000000000000",
    1953 => "000000000000000000",
    1954 => "000000000000000000",
    1955 => "000000000000000000",
    1956 => "000000000000000000",
    1957 => "000000000000000000",
    1958 => "000000000000000000",
    1959 => "000000000000000000",
    1960 => "000000000000000000",
    1961 => "000000000000000000",
    1962 => "000000000000000000",
    1963 => "000000000000000000",
    1964 => "000000000000000000",
    1965 => "000000000000000000",
    1966 => "000000000000000000",
    1967 => "000000000000000000",
    1968 => "000000000000000000",
    1969 => "000000000000000000",
    1970 => "000000000000000000",
    1971 => "000000000000000000",
    1972 => "000000000000000000",
    1973 => "000000000000000000",
    1974 => "000000000000000000",
    1975 => "000000000000000000",
    1976 => "000000000000000000",
    1977 => "000000000000000000",
    1978 => "000000000000000000",
    1979 => "000000000000000000",
    1980 => "000000000000000000",
    1981 => "000000000000000000",
    1982 => "000000000000000000",
    1983 => "000000000000000000",
    1984 => "000000000000000000",
    1985 => "000000000000000000",
    1986 => "000000000000000000",
    1987 => "000000000000000000",
    1988 => "000000000000000000",
    1989 => "000000000000000000",
    1990 => "000000000000000000",
    1991 => "000000000000000000",
    1992 => "000000000000000000",
    1993 => "000000000000000000",
    1994 => "000000000000000000",
    1995 => "000000000000000000",
    1996 => "000000000000000000",
    1997 => "000000000000000000",
    1998 => "000000000000000000",
    1999 => "000000000000000000",
    2000 => "000000000000000000",
    2001 => "000000000000000000",
    2002 => "000000000000000000",
    2003 => "000000000000000000",
    2004 => "000000000000000000",
    2005 => "000000000000000000",
    2006 => "000000000000000000",
    2007 => "000000000000000000",
    2008 => "000000000000000000",
    2009 => "000000000000000000",
    2010 => "000000000000000000",
    2011 => "000000000000000000",
    2012 => "000000000000000000",
    2013 => "000000000000000000",
    2014 => "000000000000000000",
    2015 => "000000000000000000",
    2016 => "000000000000000000",
    2017 => "000000000000000000",
    2018 => "000000000000000000",
    2019 => "000000000000000000",
    2020 => "000000000000000000",
    2021 => "000000000000000000",
    2022 => "000000000000000000",
    2023 => "000000000000000000",
    2024 => "000000000000000000",
    2025 => "000000000000000000",
    2026 => "000000000000000000",
    2027 => "000000000000000000",
    2028 => "000000000000000000",
    2029 => "000000000000000000",
    2030 => "000000000000000000",
    2031 => "000000000000000000",
    2032 => "000000000000000000",
    2033 => "000000000000000000",
    2034 => "000000000000000000",
    2035 => "000000000000000000",
    2036 => "000000000000000000",
    2037 => "000000000000000000",
    2038 => "000000000000000000",
    2039 => "000000000000000000",
    2040 => "000000000000000000",
    2041 => "000000000000000000",
    2042 => "000000000000000000",
    2043 => "000000000000000000",
    2044 => "000000000000000000",
    2045 => "000000000000000000",
    2046 => "000000000000000000",
    2047 => "000000000000000000",
    2048 => "000000000000000000",
    2049 => "000000000000000000",
    2050 => "000000000000000000",
    2051 => "000000000000000000",
    2052 => "000000000000000000",
    2053 => "000000000000000000",
    2054 => "000000000000000000",
    2055 => "000000000000000000",
    2056 => "000000000000000000",
    2057 => "000000000000000000",
    2058 => "000000000000000000",
    2059 => "000000000000000000",
    2060 => "000000000000000000",
    2061 => "000000000000000000",
    2062 => "000000000000000000",
    2063 => "000000000000000000",
    2064 => "000000000000000000",
    2065 => "000000000000000000",
    2066 => "000000000000000000",
    2067 => "000000000000000000",
    2068 => "000000000000000000",
    2069 => "000000000000000000",
    2070 => "000000000000000000",
    2071 => "000000000000000000",
    2072 => "000000000000000000",
    2073 => "000000000000000000",
    2074 => "000000000000000000",
    2075 => "000000000000000000",
    2076 => "000000000000000000",
    2077 => "000000000000000000",
    2078 => "000000000000000000",
    2079 => "000000000000000000",
    2080 => "000000000000000000",
    2081 => "000000000000000000",
    2082 => "000000000000000000",
    2083 => "000000000000000000",
    2084 => "000000000000000000",
    2085 => "000000000000000000",
    2086 => "000000000000000000",
    2087 => "000000000000000000",
    2088 => "000000000000000000",
    2089 => "000000000000000000",
    2090 => "000000000000000000",
    2091 => "000000000000000000",
    2092 => "000000000000000000",
    2093 => "000000000000000000",
    2094 => "000000000000000000",
    2095 => "000000000000000000",
    2096 => "000000000000000000",
    2097 => "000000000000000000",
    2098 => "000000000000000000",
    2099 => "000000000000000000",
    2100 => "000000000000000000",
    2101 => "000000000000000000",
    2102 => "000000000000000000",
    2103 => "000000000000000000",
    2104 => "000000000000000000",
    2105 => "000000000000000000",
    2106 => "000000000000000000",
    2107 => "000000000000000000",
    2108 => "000000000000000000",
    2109 => "000000000000000000",
    2110 => "000000000000000000",
    2111 => "000000000000000000",
    2112 => "000000000000000000",
    2113 => "000000000000000000",
    2114 => "000000000000000000",
    2115 => "000000000000000000",
    2116 => "000000000000000000",
    2117 => "000000000000000000",
    2118 => "000000000000000000",
    2119 => "000000000000000000",
    2120 => "000000000000000000",
    2121 => "000000000000000000",
    2122 => "000000000000000000",
    2123 => "000000000000000000",
    2124 => "000000000000000000",
    2125 => "000000000000000000",
    2126 => "000000000000000000",
    2127 => "000000000000000000",
    2128 => "000000000000000000",
    2129 => "000000000000000000",
    2130 => "000000000000000000",
    2131 => "000000000000000000",
    2132 => "000000000000000000",
    2133 => "000000000000000000",
    2134 => "000000000000000000",
    2135 => "000000000000000000",
    2136 => "000000000000000000",
    2137 => "000000000000000000",
    2138 => "000000000000000000",
    2139 => "000000000000000000",
    2140 => "000000000000000000",
    2141 => "000000000000000000",
    2142 => "000000000000000000",
    2143 => "000000000000000000",
    2144 => "000000000000000000",
    2145 => "000000000000000000",
    2146 => "000000000000000000",
    2147 => "000000000000000000",
    2148 => "000000000000000000",
    2149 => "000000000000000000",
    2150 => "000000000000000000",
    2151 => "000000000000000000",
    2152 => "000000000000000000",
    2153 => "000000000000000000",
    2154 => "000000000000000000",
    2155 => "000000000000000000",
    2156 => "000000000000000000",
    2157 => "000000000000000000",
    2158 => "000000000000000000",
    2159 => "000000000000000000",
    2160 => "000000000000000000",
    2161 => "000000000000000000",
    2162 => "000000000000000000",
    2163 => "000000000000000000",
    2164 => "000000000000000000",
    2165 => "000000000000000000",
    2166 => "000000000000000000",
    2167 => "000000000000000000",
    2168 => "000000000000000000",
    2169 => "000000000000000000",
    2170 => "000000000000000000",
    2171 => "000000000000000000",
    2172 => "000000000000000000",
    2173 => "000000000000000000",
    2174 => "000000000000000000",
    2175 => "000000000000000000",
    2176 => "000000000000000000",
    2177 => "000000000000000000",
    2178 => "000000000000000000",
    2179 => "000000000000000000",
    2180 => "000000000000000000",
    2181 => "000000000000000000",
    2182 => "000000000000000000",
    2183 => "000000000000000000",
    2184 => "000000000000000000",
    2185 => "000000000000000000",
    2186 => "000000000000000000",
    2187 => "000000000000000000",
    2188 => "000000000000000000",
    2189 => "000000000000000000",
    2190 => "000000000000000000",
    2191 => "000000000000000000",
    2192 => "000000000000000000",
    2193 => "000000000000000000",
    2194 => "000000000000000000",
    2195 => "000000000000000000",
    2196 => "000000000000000000",
    2197 => "000000000000000000",
    2198 => "000000000000000000",
    2199 => "000000000000000000",
    2200 => "000000000000000000",
    2201 => "000000000000000000",
    2202 => "000000000000000000",
    2203 => "000000000000000000",
    2204 => "000000000000000000",
    2205 => "000000000000000000",
    2206 => "000000000000000000",
    2207 => "000000000000000000",
    2208 => "000000000000000000",
    2209 => "000000000000000000",
    2210 => "000000000000000000",
    2211 => "000000000000000000",
    2212 => "000000000000000000",
    2213 => "000000000000000000",
    2214 => "000000000000000000",
    2215 => "000000000000000000",
    2216 => "000000000000000000",
    2217 => "000000000000000000",
    2218 => "000000000000000000",
    2219 => "000000000000000000",
    2220 => "000000000000000000",
    2221 => "000000000000000000",
    2222 => "000000000000000000",
    2223 => "000000000000000000",
    2224 => "000000000000000000",
    2225 => "000000000000000000",
    2226 => "000000000000000000",
    2227 => "000000000000000000",
    2228 => "000000000000000000",
    2229 => "000000000000000000",
    2230 => "000000000000000000",
    2231 => "000000000000000000",
    2232 => "000000000000000000",
    2233 => "000000000000000000",
    2234 => "000000000000000000",
    2235 => "000000000000000000",
    2236 => "000000000000000000",
    2237 => "000000000000000000",
    2238 => "000000000000000000",
    2239 => "000000000000000000",
    2240 => "000000000000000000",
    2241 => "000000000000000000",
    2242 => "000000000000000000",
    2243 => "000000000000000000",
    2244 => "000000000000000000",
    2245 => "000000000000000000",
    2246 => "000000000000000000",
    2247 => "000000000000000000",
    2248 => "000000000000000000",
    2249 => "000000000000000000",
    2250 => "000000000000000000",
    2251 => "000000000000000000",
    2252 => "000000000000000000",
    2253 => "000000000000000000",
    2254 => "000000000000000000",
    2255 => "000000000000000000",
    2256 => "000000000000000000",
    2257 => "000000000000000000",
    2258 => "000000000000000000",
    2259 => "000000000000000000",
    2260 => "000000000000000000",
    2261 => "000000000000000000",
    2262 => "000000000000000000",
    2263 => "000000000000000000",
    2264 => "000000000000000000",
    2265 => "000000000000000000",
    2266 => "000000000000000000",
    2267 => "000000000000000000",
    2268 => "000000000000000000",
    2269 => "000000000000000000",
    2270 => "000000000000000000",
    2271 => "000000000000000000",
    2272 => "000000000000000000",
    2273 => "000000000000000000",
    2274 => "000000000000000000",
    2275 => "000000000000000000",
    2276 => "000000000000000000",
    2277 => "000000000000000000",
    2278 => "000000000000000000",
    2279 => "000000000000000000",
    2280 => "000000000000000000",
    2281 => "000000000000000000",
    2282 => "000000000000000000",
    2283 => "000000000000000000",
    2284 => "000000000000000000",
    2285 => "000000000000000000",
    2286 => "000000000000000000",
    2287 => "000000000000000000",
    2288 => "000000000000000000",
    2289 => "000000000000000000",
    2290 => "000000000000000000",
    2291 => "000000000000000000",
    2292 => "000000000000000000",
    2293 => "000000000000000000",
    2294 => "000000000000000000",
    2295 => "000000000000000000",
    2296 => "000000000000000000",
    2297 => "000000000000000000",
    2298 => "000000000000000000",
    2299 => "000000000000000000",
    2300 => "000000000000000000",
    2301 => "000000000000000000",
    2302 => "000000000000000000",
    2303 => "000000000000000000",
    2304 => "000000000000000000",
    2305 => "000000000000000000",
    2306 => "000000000000000000",
    2307 => "000000000000000000",
    2308 => "000000000000000000",
    2309 => "000000000000000000",
    2310 => "000000000000000000",
    2311 => "000000000000000000",
    2312 => "000000000000000000",
    2313 => "000000000000000000",
    2314 => "000000000000000000",
    2315 => "000000000000000000",
    2316 => "000000000000000000",
    2317 => "000000000000000000",
    2318 => "000000000000000000",
    2319 => "000000000000000000",
    2320 => "000000000000000000",
    2321 => "000000000000000000",
    2322 => "000000000000000000",
    2323 => "000000000000000000",
    2324 => "000000000000000000",
    2325 => "000000000000000000",
    2326 => "000000000000000000",
    2327 => "000000000000000000",
    2328 => "000000000000000000",
    2329 => "000000000000000000",
    2330 => "000000000000000000",
    2331 => "000000000000000000",
    2332 => "000000000000000000",
    2333 => "000000000000000000",
    2334 => "000000000000000000",
    2335 => "000000000000000000",
    2336 => "000000000000000000",
    2337 => "000000000000000000",
    2338 => "000000000000000000",
    2339 => "000000000000000000",
    2340 => "000000000000000000",
    2341 => "000000000000000000",
    2342 => "000000000000000000",
    2343 => "000000000000000000",
    2344 => "000000000000000000",
    2345 => "000000000000000000",
    2346 => "000000000000000000",
    2347 => "000000000000000000",
    2348 => "000000000000000000",
    2349 => "000000000000000000",
    2350 => "000000000000000000",
    2351 => "000000000000000000",
    2352 => "000000000000000000",
    2353 => "000000000000000000",
    2354 => "000000000000000000",
    2355 => "000000000000000000",
    2356 => "000000000000000000",
    2357 => "000000000000000000",
    2358 => "000000000000000000",
    2359 => "000000000000000000",
    2360 => "000000000000000000",
    2361 => "000000000000000000",
    2362 => "000000000000000000",
    2363 => "000000000000000000",
    2364 => "000000000000000000",
    2365 => "000000000000000000",
    2366 => "000000000000000000",
    2367 => "000000000000000000",
    2368 => "000000000000000000",
    2369 => "000000000000000000",
    2370 => "000000000000000000",
    2371 => "000000000000000000",
    2372 => "000000000000000000",
    2373 => "000000000000000000",
    2374 => "000000000000000000",
    2375 => "000000000000000000",
    2376 => "000000000000000000",
    2377 => "000000000000000000",
    2378 => "000000000000000000",
    2379 => "000000000000000000",
    2380 => "000000000000000000",
    2381 => "000000000000000000",
    2382 => "000000000000000000",
    2383 => "000000000000000000",
    2384 => "000000000000000000",
    2385 => "000000000000000000",
    2386 => "000000000000000000",
    2387 => "000000000000000000",
    2388 => "000000000000000000",
    2389 => "000000000000000000",
    2390 => "000000000000000000",
    2391 => "000000000000000000",
    2392 => "000000000000000000",
    2393 => "000000000000000000",
    2394 => "000000000000000000",
    2395 => "000000000000000000",
    2396 => "000000000000000000",
    2397 => "000000000000000000",
    2398 => "000000000000000000",
    2399 => "000000000000000000",
    2400 => "000000000000000000",
    2401 => "000000000000000000",
    2402 => "000000000000000000",
    2403 => "000000000000000000",
    2404 => "000000000000000000",
    2405 => "000000000000000000",
    2406 => "000000000000000000",
    2407 => "000000000000000000",
    2408 => "000000000000000000",
    2409 => "000000000000000000",
    2410 => "000000000000000000",
    2411 => "000000000000000000",
    2412 => "000000000000000000",
    2413 => "000000000000000000",
    2414 => "000000000000000000",
    2415 => "000000000000000000",
    2416 => "000000000000000000",
    2417 => "000000000000000000",
    2418 => "000000000000000000",
    2419 => "000000000000000000",
    2420 => "000000000000000000",
    2421 => "000000000000000000",
    2422 => "000000000000000000",
    2423 => "000000000000000000",
    2424 => "000000000000000000",
    2425 => "000000000000000000",
    2426 => "000000000000000000",
    2427 => "000000000000000000",
    2428 => "000000000000000000",
    2429 => "000000000000000000",
    2430 => "000000000000000000",
    2431 => "000000000000000000",
    2432 => "000000000000000000",
    2433 => "000000000000000000",
    2434 => "000000000000000000",
    2435 => "000000000000000000",
    2436 => "000000000000000000",
    2437 => "000000000000000000",
    2438 => "000000000000000000",
    2439 => "000000000000000000",
    2440 => "000000000000000000",
    2441 => "000000000000000000",
    2442 => "000000000000000000",
    2443 => "000000000000000000",
    2444 => "000000000000000000",
    2445 => "000000000000000000",
    2446 => "000000000000000000",
    2447 => "000000000000000000",
    2448 => "000000000000000000",
    2449 => "000000000000000000",
    2450 => "000000000000000000",
    2451 => "000000000000000000",
    2452 => "000000000000000000",
    2453 => "000000000000000000",
    2454 => "000000000000000000",
    2455 => "000000000000000000",
    2456 => "000000000000000000",
    2457 => "000000000000000000",
    2458 => "000000000000000000",
    2459 => "000000000000000000",
    2460 => "000000000000000000",
    2461 => "000000000000000000",
    2462 => "000000000000000000",
    2463 => "000000000000000000",
    2464 => "000000000000000000",
    2465 => "000000000000000000",
    2466 => "000000000000000000",
    2467 => "000000000000000000",
    2468 => "000000000000000000",
    2469 => "000000000000000000",
    2470 => "000000000000000000",
    2471 => "000000000000000000",
    2472 => "000000000000000000",
    2473 => "000000000000000000",
    2474 => "000000000000000000",
    2475 => "000000000000000000",
    2476 => "000000000000000000",
    2477 => "000000000000000000",
    2478 => "000000000000000000",
    2479 => "000000000000000000",
    2480 => "000000000000000000",
    2481 => "000000000000000000",
    2482 => "000000000000000000",
    2483 => "000000000000000000",
    2484 => "000000000000000000",
    2485 => "000000000000000000",
    2486 => "000000000000000000",
    2487 => "000000000000000000",
    2488 => "000000000000000000",
    2489 => "000000000000000000",
    2490 => "000000000000000000",
    2491 => "000000000000000000",
    2492 => "000000000000000000",
    2493 => "000000000000000000",
    2494 => "000000000000000000",
    2495 => "000000000000000000",
    2496 => "000000000000000000",
    2497 => "000000000000000000",
    2498 => "000000000000000000",
    2499 => "000000000000000000",
    2500 => "000000000000000000",
    2501 => "000000000000000000",
    2502 => "000000000000000000",
    2503 => "000000000000000000",
    2504 => "000000000000000000",
    2505 => "000000000000000000",
    2506 => "000000000000000000",
    2507 => "000000000000000000",
    2508 => "000000000000000000",
    2509 => "000000000000000000",
    2510 => "000000000000000000",
    2511 => "000000000000000000",
    2512 => "000000000000000000",
    2513 => "000000000000000000",
    2514 => "000000000000000000",
    2515 => "000000000000000000",
    2516 => "000000000000000000",
    2517 => "000000000000000000",
    2518 => "000000000000000000",
    2519 => "000000000000000000",
    2520 => "000000000000000000",
    2521 => "000000000000000000",
    2522 => "000000000000000000",
    2523 => "000000000000000000",
    2524 => "000000000000000000",
    2525 => "000000000000000000",
    2526 => "000000000000000000",
    2527 => "000000000000000000",
    2528 => "000000000000000000",
    2529 => "000000000000000000",
    2530 => "000000000000000000",
    2531 => "000000000000000000",
    2532 => "000000000000000000",
    2533 => "000000000000000000",
    2534 => "000000000000000000",
    2535 => "000000000000000000",
    2536 => "000000000000000000",
    2537 => "000000000000000000",
    2538 => "000000000000000000",
    2539 => "000000000000000000",
    2540 => "000000000000000000",
    2541 => "000000000000000000",
    2542 => "000000000000000000",
    2543 => "000000000000000000",
    2544 => "000000000000000000",
    2545 => "000000000000000000",
    2546 => "000000000000000000",
    2547 => "000000000000000000",
    2548 => "000000000000000000",
    2549 => "000000000000000000",
    2550 => "000000000000000000",
    2551 => "000000000000000000",
    2552 => "000000000000000000",
    2553 => "000000000000000000",
    2554 => "000000000000000000",
    2555 => "000000000000000000",
    2556 => "000000000000000000",
    2557 => "000000000000000000",
    2558 => "000000000000000000",
    2559 => "000000000000000000",
    2560 => "000000000000000000",
    2561 => "000000000000000000",
    2562 => "000000000000000000",
    2563 => "000000000000000000",
    2564 => "000000000000000000",
    2565 => "000000000000000000",
    2566 => "000000000000000000",
    2567 => "000000000000000000",
    2568 => "000000000000000000",
    2569 => "000000000000000000",
    2570 => "000000000000000000",
    2571 => "000000000000000000",
    2572 => "000000000000000000",
    2573 => "000000000000000000",
    2574 => "000000000000000000",
    2575 => "000000000000000000",
    2576 => "000000000000000000",
    2577 => "000000000000000000",
    2578 => "000000000000000000",
    2579 => "000000000000000000",
    2580 => "000000000000000000",
    2581 => "000000000000000000",
    2582 => "000000000000000000",
    2583 => "000000000000000000",
    2584 => "000000000000000000",
    2585 => "000000000000000000",
    2586 => "000000000000000000",
    2587 => "000000000000000000",
    2588 => "000000000000000000",
    2589 => "000000000000000000",
    2590 => "000000000000000000",
    2591 => "000000000000000000",
    2592 => "000000000000000000",
    2593 => "000000000000000000",
    2594 => "000000000000000000",
    2595 => "000000000000000000",
    2596 => "000000000000000000",
    2597 => "000000000000000000",
    2598 => "000000000000000000",
    2599 => "000000000000000000",
    2600 => "000000000000000000",
    2601 => "000000000000000000",
    2602 => "000000000000000000",
    2603 => "000000000000000000",
    2604 => "000000000000000000",
    2605 => "000000000000000000",
    2606 => "000000000000000000",
    2607 => "000000000000000000",
    2608 => "000000000000000000",
    2609 => "000000000000000000",
    2610 => "000000000000000000",
    2611 => "000000000000000000",
    2612 => "000000000000000000",
    2613 => "000000000000000000",
    2614 => "000000000000000000",
    2615 => "000000000000000000",
    2616 => "000000000000000000",
    2617 => "000000000000000000",
    2618 => "000000000000000000",
    2619 => "000000000000000000",
    2620 => "000000000000000000",
    2621 => "000000000000000000",
    2622 => "000000000000000000",
    2623 => "000000000000000000",
    2624 => "000000000000000000",
    2625 => "000000000000000000",
    2626 => "000000000000000000",
    2627 => "000000000000000000",
    2628 => "000000000000000000",
    2629 => "000000000000000000",
    2630 => "000000000000000000",
    2631 => "000000000000000000",
    2632 => "000000000000000000",
    2633 => "000000000000000000",
    2634 => "000000000000000000",
    2635 => "000000000000000000",
    2636 => "000000000000000000",
    2637 => "000000000000000000",
    2638 => "000000000000000000",
    2639 => "000000000000000000",
    2640 => "000000000000000000",
    2641 => "000000000000000000",
    2642 => "000000000000000000",
    2643 => "000000000000000000",
    2644 => "000000000000000000",
    2645 => "000000000000000000",
    2646 => "000000000000000000",
    2647 => "000000000000000000",
    2648 => "000000000000000000",
    2649 => "000000000000000000",
    2650 => "000000000000000000",
    2651 => "000000000000000000",
    2652 => "000000000000000000",
    2653 => "000000000000000000",
    2654 => "000000000000000000",
    2655 => "000000000000000000",
    2656 => "000000000000000000",
    2657 => "000000000000000000",
    2658 => "000000000000000000",
    2659 => "000000000000000000",
    2660 => "000000000000000000",
    2661 => "000000000000000000",
    2662 => "000000000000000000",
    2663 => "000000000000000000",
    2664 => "000000000000000000",
    2665 => "000000000000000000",
    2666 => "000000000000000000",
    2667 => "000000000000000000",
    2668 => "000000000000000000",
    2669 => "000000000000000000",
    2670 => "000000000000000000",
    2671 => "000000000000000000",
    2672 => "000000000000000000",
    2673 => "000000000000000000",
    2674 => "000000000000000000",
    2675 => "000000000000000000",
    2676 => "000000000000000000",
    2677 => "000000000000000000",
    2678 => "000000000000000000",
    2679 => "000000000000000000",
    2680 => "000000000000000000",
    2681 => "000000000000000000",
    2682 => "000000000000000000",
    2683 => "000000000000000000",
    2684 => "000000000000000000",
    2685 => "000000000000000000",
    2686 => "000000000000000000",
    2687 => "000000000000000000",
    2688 => "000000000000000000",
    2689 => "000000000000000000",
    2690 => "000000000000000000",
    2691 => "000000000000000000",
    2692 => "000000000000000000",
    2693 => "000000000000000000",
    2694 => "000000000000000000",
    2695 => "000000000000000000",
    2696 => "000000000000000000",
    2697 => "000000000000000000",
    2698 => "000000000000000000",
    2699 => "000000000000000000",
    2700 => "000000000000000000",
    2701 => "000000000000000000",
    2702 => "000000000000000000",
    2703 => "000000000000000000",
    2704 => "000000000000000000",
    2705 => "000000000000000000",
    2706 => "000000000000000000",
    2707 => "000000000000000000",
    2708 => "000000000000000000",
    2709 => "000000000000000000",
    2710 => "000000000000000000",
    2711 => "000000000000000000",
    2712 => "000000000000000000",
    2713 => "000000000000000000",
    2714 => "000000000000000000",
    2715 => "000000000000000000",
    2716 => "000000000000000000",
    2717 => "000000000000000000",
    2718 => "000000000000000000",
    2719 => "000000000000000000",
    2720 => "000000000000000000",
    2721 => "000000000000000000",
    2722 => "000000000000000000",
    2723 => "000000000000000000",
    2724 => "000000000000000000",
    2725 => "000000000000000000",
    2726 => "000000000000000000",
    2727 => "000000000000000000",
    2728 => "000000000000000000",
    2729 => "000000000000000000",
    2730 => "000000000000000000",
    2731 => "000000000000000000",
    2732 => "000000000000000000",
    2733 => "000000000000000000",
    2734 => "000000000000000000",
    2735 => "000000000000000000",
    2736 => "000000000000000000",
    2737 => "000000000000000000",
    2738 => "000000000000000000",
    2739 => "000000000000000000",
    2740 => "000000000000000000",
    2741 => "000000000000000000",
    2742 => "000000000000000000",
    2743 => "000000000000000000",
    2744 => "000000000000000000",
    2745 => "000000000000000000",
    2746 => "000000000000000000",
    2747 => "000000000000000000",
    2748 => "000000000000000000",
    2749 => "000000000000000000",
    2750 => "000000000000000000",
    2751 => "000000000000000000",
    2752 => "000000000000000000",
    2753 => "000000000000000000",
    2754 => "000000000000000000",
    2755 => "000000000000000000",
    2756 => "000000000000000000",
    2757 => "000000000000000000",
    2758 => "000000000000000000",
    2759 => "000000000000000000",
    2760 => "000000000000000000",
    2761 => "000000000000000000",
    2762 => "000000000000000000",
    2763 => "000000000000000000",
    2764 => "000000000000000000",
    2765 => "000000000000000000",
    2766 => "000000000000000000",
    2767 => "000000000000000000",
    2768 => "000000000000000000",
    2769 => "000000000000000000",
    2770 => "000000000000000000",
    2771 => "000000000000000000",
    2772 => "000000000000000000",
    2773 => "000000000000000000",
    2774 => "000000000000000000",
    2775 => "000000000000000000",
    2776 => "000000000000000000",
    2777 => "000000000000000000",
    2778 => "000000000000000000",
    2779 => "000000000000000000",
    2780 => "000000000000000000",
    2781 => "000000000000000000",
    2782 => "000000000000000000",
    2783 => "000000000000000000",
    2784 => "000000000000000000",
    2785 => "000000000000000000",
    2786 => "000000000000000000",
    2787 => "000000000000000000",
    2788 => "000000000000000000",
    2789 => "000000000000000000",
    2790 => "000000000000000000",
    2791 => "000000000000000000",
    2792 => "000000000000000000",
    2793 => "000000000000000000",
    2794 => "000000000000000000",
    2795 => "000000000000000000",
    2796 => "000000000000000000",
    2797 => "000000000000000000",
    2798 => "000000000000000000",
    2799 => "000000000000000000",
    2800 => "000000000000000000",
    2801 => "000000000000000000",
    2802 => "000000000000000000",
    2803 => "000000000000000000",
    2804 => "000000000000000000",
    2805 => "000000000000000000",
    2806 => "000000000000000000",
    2807 => "000000000000000000",
    2808 => "000000000000000000",
    2809 => "000000000000000000",
    2810 => "000000000000000000",
    2811 => "000000000000000000",
    2812 => "000000000000000000",
    2813 => "000000000000000000",
    2814 => "000000000000000000",
    2815 => "000000000000000000",
    2816 => "000000000000000000",
    2817 => "000000000000000000",
    2818 => "000000000000000000",
    2819 => "000000000000000000",
    2820 => "000000000000000000",
    2821 => "000000000000000000",
    2822 => "000000000000000000",
    2823 => "000000000000000000",
    2824 => "000000000000000000",
    2825 => "000000000000000000",
    2826 => "000000000000000000",
    2827 => "000000000000000000",
    2828 => "000000000000000000",
    2829 => "000000000000000000",
    2830 => "000000000000000000",
    2831 => "000000000000000000",
    2832 => "000000000000000000",
    2833 => "000000000000000000",
    2834 => "000000000000000000",
    2835 => "000000000000000000",
    2836 => "000000000000000000",
    2837 => "000000000000000000",
    2838 => "000000000000000000",
    2839 => "000000000000000000",
    2840 => "000000000000000000",
    2841 => "000000000000000000",
    2842 => "000000000000000000",
    2843 => "000000000000000000",
    2844 => "000000000000000000",
    2845 => "000000000000000000",
    2846 => "000000000000000000",
    2847 => "000000000000000000",
    2848 => "000000000000000000",
    2849 => "000000000000000000",
    2850 => "000000000000000000",
    2851 => "000000000000000000",
    2852 => "000000000000000000",
    2853 => "000000000000000000",
    2854 => "000000000000000000",
    2855 => "000000000000000000",
    2856 => "000000000000000000",
    2857 => "000000000000000000",
    2858 => "000000000000000000",
    2859 => "000000000000000000",
    2860 => "000000000000000000",
    2861 => "000000000000000000",
    2862 => "000000000000000000",
    2863 => "000000000000000000",
    2864 => "000000000000000000",
    2865 => "000000000000000000",
    2866 => "000000000000000000",
    2867 => "000000000000000000",
    2868 => "000000000000000000",
    2869 => "000000000000000000",
    2870 => "000000000000000000",
    2871 => "000000000000000000",
    2872 => "000000000000000000",
    2873 => "000000000000000000",
    2874 => "000000000000000000",
    2875 => "000000000000000000",
    2876 => "000000000000000000",
    2877 => "000000000000000000",
    2878 => "000000000000000000",
    2879 => "000000000000000000",
    2880 => "000000000000000000",
    2881 => "000000000000000000",
    2882 => "000000000000000000",
    2883 => "000000000000000000",
    2884 => "000000000000000000",
    2885 => "000000000000000000",
    2886 => "000000000000000000",
    2887 => "000000000000000000",
    2888 => "000000000000000000",
    2889 => "000000000000000000",
    2890 => "000000000000000000",
    2891 => "000000000000000000",
    2892 => "000000000000000000",
    2893 => "000000000000000000",
    2894 => "000000000000000000",
    2895 => "000000000000000000",
    2896 => "000000000000000000",
    2897 => "000000000000000000",
    2898 => "000000000000000000",
    2899 => "000000000000000000",
    2900 => "000000000000000000",
    2901 => "000000000000000000",
    2902 => "000000000000000000",
    2903 => "000000000000000000",
    2904 => "000000000000000000",
    2905 => "000000000000000000",
    2906 => "000000000000000000",
    2907 => "000000000000000000",
    2908 => "000000000000000000",
    2909 => "000000000000000000",
    2910 => "000000000000000000",
    2911 => "000000000000000000",
    2912 => "000000000000000000",
    2913 => "000000000000000000",
    2914 => "000000000000000000",
    2915 => "000000000000000000",
    2916 => "000000000000000000",
    2917 => "000000000000000000",
    2918 => "000000000000000000",
    2919 => "000000000000000000",
    2920 => "000000000000000000",
    2921 => "000000000000000000",
    2922 => "000000000000000000",
    2923 => "000000000000000000",
    2924 => "000000000000000000",
    2925 => "000000000000000000",
    2926 => "000000000000000000",
    2927 => "000000000000000000",
    2928 => "000000000000000000",
    2929 => "000000000000000000",
    2930 => "000000000000000000",
    2931 => "000000000000000000",
    2932 => "000000000000000000",
    2933 => "000000000000000000",
    2934 => "000000000000000000",
    2935 => "000000000000000000",
    2936 => "000000000000000000",
    2937 => "000000000000000000",
    2938 => "000000000000000000",
    2939 => "000000000000000000",
    2940 => "000000000000000000",
    2941 => "000000000000000000",
    2942 => "000000000000000000",
    2943 => "000000000000000000",
    2944 => "000000000000000000",
    2945 => "000000000000000000",
    2946 => "000000000000000000",
    2947 => "000000000000000000",
    2948 => "000000000000000000",
    2949 => "000000000000000000",
    2950 => "000000000000000000",
    2951 => "000000000000000000",
    2952 => "000000000000000000",
    2953 => "000000000000000000",
    2954 => "000000000000000000",
    2955 => "000000000000000000",
    2956 => "000000000000000000",
    2957 => "000000000000000000",
    2958 => "000000000000000000",
    2959 => "000000000000000000",
    2960 => "000000000000000000",
    2961 => "000000000000000000",
    2962 => "000000000000000000",
    2963 => "000000000000000000",
    2964 => "000000000000000000",
    2965 => "000000000000000000",
    2966 => "000000000000000000",
    2967 => "000000000000000000",
    2968 => "000000000000000000",
    2969 => "000000000000000000",
    2970 => "000000000000000000",
    2971 => "000000000000000000",
    2972 => "000000000000000000",
    2973 => "000000000000000000",
    2974 => "000000000000000000",
    2975 => "000000000000000000",
    2976 => "000000000000000000",
    2977 => "000000000000000000",
    2978 => "000000000000000000",
    2979 => "000000000000000000",
    2980 => "000000000000000000",
    2981 => "000000000000000000",
    2982 => "000000000000000000",
    2983 => "000000000000000000",
    2984 => "000000000000000000",
    2985 => "000000000000000000",
    2986 => "000000000000000000",
    2987 => "000000000000000000",
    2988 => "000000000000000000",
    2989 => "000000000000000000",
    2990 => "000000000000000000",
    2991 => "000000000000000000",
    2992 => "000000000000000000",
    2993 => "000000000000000000",
    2994 => "000000000000000000",
    2995 => "000000000000000000",
    2996 => "000000000000000000",
    2997 => "000000000000000000",
    2998 => "000000000000000000",
    2999 => "000000000000000000",
    3000 => "000000000000000000",
    3001 => "000000000000000000",
    3002 => "000000000000000000",
    3003 => "000000000000000000",
    3004 => "000000000000000000",
    3005 => "000000000000000000",
    3006 => "000000000000000000",
    3007 => "000000000000000000",
    3008 => "000000000000000000",
    3009 => "000000000000000000",
    3010 => "000000000000000000",
    3011 => "000000000000000000",
    3012 => "000000000000000000",
    3013 => "000000000000000000",
    3014 => "000000000000000000",
    3015 => "000000000000000000",
    3016 => "000000000000000000",
    3017 => "000000000000000000",
    3018 => "000000000000000000",
    3019 => "000000000000000000",
    3020 => "000000000000000000",
    3021 => "000000000000000000",
    3022 => "000000000000000000",
    3023 => "000000000000000000",
    3024 => "000000000000000000",
    3025 => "000000000000000000",
    3026 => "000000000000000000",
    3027 => "000000000000000000",
    3028 => "000000000000000000",
    3029 => "000000000000000000",
    3030 => "000000000000000000",
    3031 => "000000000000000000",
    3032 => "000000000000000000",
    3033 => "000000000000000000",
    3034 => "000000000000000000",
    3035 => "000000000000000000",
    3036 => "000000000000000000",
    3037 => "000000000000000000",
    3038 => "000000000000000000",
    3039 => "000000000000000000",
    3040 => "000000000000000000",
    3041 => "000000000000000000",
    3042 => "000000000000000000",
    3043 => "000000000000000000",
    3044 => "000000000000000000",
    3045 => "000000000000000000",
    3046 => "000000000000000000",
    3047 => "000000000000000000",
    3048 => "000000000000000000",
    3049 => "000000000000000000",
    3050 => "000000000000000000",
    3051 => "000000000000000000",
    3052 => "000000000000000000",
    3053 => "000000000000000000",
    3054 => "000000000000000000",
    3055 => "000000000000000000",
    3056 => "000000000000000000",
    3057 => "000000000000000000",
    3058 => "000000000000000000",
    3059 => "000000000000000000",
    3060 => "000000000000000000",
    3061 => "000000000000000000",
    3062 => "000000000000000000",
    3063 => "000000000000000000",
    3064 => "000000000000000000",
    3065 => "000000000000000000",
    3066 => "000000000000000000",
    3067 => "000000000000000000",
    3068 => "000000000000000000",
    3069 => "000000000000000000",
    3070 => "000000000000000000",
    3071 => "000000000000000000",
    3072 => "000000000000000000",
    3073 => "000000000000000000",
    3074 => "000000000000000000",
    3075 => "000000000000000000",
    3076 => "000000000000000000",
    3077 => "000000000000000000",
    3078 => "000000000000000000",
    3079 => "000000000000000000",
    3080 => "000000000000000000",
    3081 => "000000000000000000",
    3082 => "000000000000000000",
    3083 => "000000000000000000",
    3084 => "000000000000000000",
    3085 => "000000000000000000",
    3086 => "000000000000000000",
    3087 => "000000000000000000",
    3088 => "000000000000000000",
    3089 => "000000000000000000",
    3090 => "000000000000000000",
    3091 => "000000000000000000",
    3092 => "000000000000000000",
    3093 => "000000000000000000",
    3094 => "000000000000000000",
    3095 => "000000000000000000",
    3096 => "000000000000000000",
    3097 => "000000000000000000",
    3098 => "000000000000000000",
    3099 => "000000000000000000",
    3100 => "000000000000000000",
    3101 => "000000000000000000",
    3102 => "000000000000000000",
    3103 => "000000000000000000",
    3104 => "000000000000000000",
    3105 => "000000000000000000",
    3106 => "000000000000000000",
    3107 => "000000000000000000",
    3108 => "000000000000000000",
    3109 => "000000000000000000",
    3110 => "000000000000000000",
    3111 => "000000000000000000",
    3112 => "000000000000000000",
    3113 => "000000000000000000",
    3114 => "000000000000000000",
    3115 => "000000000000000000",
    3116 => "000000000000000000",
    3117 => "000000000000000000",
    3118 => "000000000000000000",
    3119 => "000000000000000000",
    3120 => "000000000000000000",
    3121 => "000000000000000000",
    3122 => "000000000000000000",
    3123 => "000000000000000000",
    3124 => "000000000000000000",
    3125 => "000000000000000000",
    3126 => "000000000000000000",
    3127 => "000000000000000000",
    3128 => "000000000000000000",
    3129 => "000000000000000000",
    3130 => "000000000000000000",
    3131 => "000000000000000000",
    3132 => "000000000000000000",
    3133 => "000000000000000000",
    3134 => "000000000000000000",
    3135 => "000000000000000000",
    3136 => "000000000000000000",
    3137 => "000000000000000000",
    3138 => "000000000000000000",
    3139 => "000000000000000000",
    3140 => "000000000000000000",
    3141 => "000000000000000000",
    3142 => "000000000000000000",
    3143 => "000000000000000000",
    3144 => "000000000000000000",
    3145 => "000000000000000000",
    3146 => "000000000000000000",
    3147 => "000000000000000000",
    3148 => "000000000000000000",
    3149 => "000000000000000000",
    3150 => "000000000000000000",
    3151 => "000000000000000000",
    3152 => "000000000000000000",
    3153 => "000000000000000000",
    3154 => "000000000000000000",
    3155 => "000000000000000000",
    3156 => "000000000000000000",
    3157 => "000000000000000000",
    3158 => "000000000000000000",
    3159 => "000000000000000000",
    3160 => "000000000000000000",
    3161 => "000000000000000000",
    3162 => "000000000000000000",
    3163 => "000000000000000000",
    3164 => "000000000000000000",
    3165 => "000000000000000000",
    3166 => "000000000000000000",
    3167 => "000000000000000000",
    3168 => "000000000000000000",
    3169 => "000000000000000000",
    3170 => "000000000000000000",
    3171 => "000000000000000000",
    3172 => "000000000000000000",
    3173 => "000000000000000000",
    3174 => "000000000000000000",
    3175 => "000000000000000000",
    3176 => "000000000000000000",
    3177 => "000000000000000000",
    3178 => "000000000000000000",
    3179 => "000000000000000000",
    3180 => "000000000000000000",
    3181 => "000000000000000000",
    3182 => "000000000000000000",
    3183 => "000000000000000000",
    3184 => "000000000000000000",
    3185 => "000000000000000000",
    3186 => "000000000000000000",
    3187 => "000000000000000000",
    3188 => "000000000000000000",
    3189 => "000000000000000000",
    3190 => "000000000000000000",
    3191 => "000000000000000000",
    3192 => "000000000000000000",
    3193 => "000000000000000000",
    3194 => "000000000000000000",
    3195 => "000000000000000000",
    3196 => "000000000000000000",
    3197 => "000000000000000000",
    3198 => "000000000000000000",
    3199 => "000000000000000000",
    3200 => "000000000000000000",
    3201 => "000000000000000000",
    3202 => "000000000000000000",
    3203 => "000000000000000000",
    3204 => "000000000000000000",
    3205 => "000000000000000000",
    3206 => "000000000000000000",
    3207 => "000000000000000000",
    3208 => "000000000000000000",
    3209 => "000000000000000000",
    3210 => "000000000000000000",
    3211 => "000000000000000000",
    3212 => "000000000000000000",
    3213 => "000000000000000000",
    3214 => "000000000000000000",
    3215 => "000000000000000000",
    3216 => "000000000000000000",
    3217 => "000000000000000000",
    3218 => "000000000000000000",
    3219 => "000000000000000000",
    3220 => "000000000000000000",
    3221 => "000000000000000000",
    3222 => "000000000000000000",
    3223 => "000000000000000000",
    3224 => "000000000000000000",
    3225 => "000000000000000000",
    3226 => "000000000000000000",
    3227 => "000000000000000000",
    3228 => "000000000000000000",
    3229 => "000000000000000000",
    3230 => "000000000000000000",
    3231 => "000000000000000000",
    3232 => "000000000000000000",
    3233 => "000000000000000000",
    3234 => "000000000000000000",
    3235 => "000000000000000000",
    3236 => "000000000000000000",
    3237 => "000000000000000000",
    3238 => "000000000000000000",
    3239 => "000000000000000000",
    3240 => "000000000000000000",
    3241 => "000000000000000000",
    3242 => "000000000000000000",
    3243 => "000000000000000000",
    3244 => "000000000000000000",
    3245 => "000000000000000000",
    3246 => "000000000000000000",
    3247 => "000000000000000000",
    3248 => "000000000000000000",
    3249 => "000000000000000000",
    3250 => "000000000000000000",
    3251 => "000000000000000000",
    3252 => "000000000000000000",
    3253 => "000000000000000000",
    3254 => "000000000000000000",
    3255 => "000000000000000000",
    3256 => "000000000000000000",
    3257 => "000000000000000000",
    3258 => "000000000000000000",
    3259 => "000000000000000000",
    3260 => "000000000000000000",
    3261 => "000000000000000000",
    3262 => "000000000000000000",
    3263 => "000000000000000000",
    3264 => "000000000000000000",
    3265 => "000000000000000000",
    3266 => "000000000000000000",
    3267 => "000000000000000000",
    3268 => "000000000000000000",
    3269 => "000000000000000000",
    3270 => "000000000000000000",
    3271 => "000000000000000000",
    3272 => "000000000000000000",
    3273 => "000000000000000000",
    3274 => "000000000000000000",
    3275 => "000000000000000000",
    3276 => "000000000000000000",
    3277 => "000000000000000000",
    3278 => "000000000000000000",
    3279 => "000000000000000000",
    3280 => "000000000000000000",
    3281 => "000000000000000000",
    3282 => "000000000000000000",
    3283 => "000000000000000000",
    3284 => "000000000000000000",
    3285 => "000000000000000000",
    3286 => "000000000000000000",
    3287 => "000000000000000000",
    3288 => "000000000000000000",
    3289 => "000000000000000000",
    3290 => "000000000000000000",
    3291 => "000000000000000000",
    3292 => "000000000000000000",
    3293 => "000000000000000000",
    3294 => "000000000000000000",
    3295 => "000000000000000000",
    3296 => "000000000000000000",
    3297 => "000000000000000000",
    3298 => "000000000000000000",
    3299 => "000000000000000000",
    3300 => "000000000000000000",
    3301 => "000000000000000000",
    3302 => "000000000000000000",
    3303 => "000000000000000000",
    3304 => "000000000000000000",
    3305 => "000000000000000000",
    3306 => "000000000000000000",
    3307 => "000000000000000000",
    3308 => "000000000000000000",
    3309 => "000000000000000000",
    3310 => "000000000000000000",
    3311 => "000000000000000000",
    3312 => "000000000000000000",
    3313 => "000000000000000000",
    3314 => "000000000000000000",
    3315 => "000000000000000000",
    3316 => "000000000000000000",
    3317 => "000000000000000000",
    3318 => "000000000000000000",
    3319 => "000000000000000000",
    3320 => "000000000000000000",
    3321 => "000000000000000000",
    3322 => "000000000000000000",
    3323 => "000000000000000000",
    3324 => "000000000000000000",
    3325 => "000000000000000000",
    3326 => "000000000000000000",
    3327 => "000000000000000000",
    3328 => "000000000000000000",
    3329 => "000000000000000000",
    3330 => "000000000000000000",
    3331 => "000000000000000000",
    3332 => "000000000000000000",
    3333 => "000000000000000000",
    3334 => "000000000000000000",
    3335 => "000000000000000000",
    3336 => "000000000000000000",
    3337 => "000000000000000000",
    3338 => "000000000000000000",
    3339 => "000000000000000000",
    3340 => "000000000000000000",
    3341 => "000000000000000000",
    3342 => "000000000000000000",
    3343 => "000000000000000000",
    3344 => "000000000000000000",
    3345 => "000000000000000000",
    3346 => "000000000000000000",
    3347 => "000000000000000000",
    3348 => "000000000000000000",
    3349 => "000000000000000000",
    3350 => "000000000000000000",
    3351 => "000000000000000000",
    3352 => "000000000000000000",
    3353 => "000000000000000000",
    3354 => "000000000000000000",
    3355 => "000000000000000000",
    3356 => "000000000000000000",
    3357 => "000000000000000000",
    3358 => "000000000000000000",
    3359 => "000000000000000000",
    3360 => "000000000000000000",
    3361 => "000000000000000000",
    3362 => "000000000000000000",
    3363 => "000000000000000000",
    3364 => "000000000000000000",
    3365 => "000000000000000000",
    3366 => "000000000000000000",
    3367 => "000000000000000000",
    3368 => "000000000000000000",
    3369 => "000000000000000000",
    3370 => "000000000000000000",
    3371 => "000000000000000000",
    3372 => "000000000000000000",
    3373 => "000000000000000000",
    3374 => "000000000000000000",
    3375 => "000000000000000000",
    3376 => "000000000000000000",
    3377 => "000000000000000000",
    3378 => "000000000000000000",
    3379 => "000000000000000000",
    3380 => "000000000000000000",
    3381 => "000000000000000000",
    3382 => "000000000000000000",
    3383 => "000000000000000000",
    3384 => "000000000000000000",
    3385 => "000000000000000000",
    3386 => "000000000000000000",
    3387 => "000000000000000000",
    3388 => "000000000000000000",
    3389 => "000000000000000000",
    3390 => "000000000000000000",
    3391 => "000000000000000000",
    3392 => "000000000000000000",
    3393 => "000000000000000000",
    3394 => "000000000000000000",
    3395 => "000000000000000000",
    3396 => "000000000000000000",
    3397 => "000000000000000000",
    3398 => "000000000000000000",
    3399 => "000000000000000000",
    3400 => "000000000000000000",
    3401 => "000000000000000000",
    3402 => "000000000000000000",
    3403 => "000000000000000000",
    3404 => "000000000000000000",
    3405 => "000000000000000000",
    3406 => "000000000000000000",
    3407 => "000000000000000000",
    3408 => "000000000000000000",
    3409 => "000000000000000000",
    3410 => "000000000000000000",
    3411 => "000000000000000000",
    3412 => "000000000000000000",
    3413 => "000000000000000000",
    3414 => "000000000000000000",
    3415 => "000000000000000000",
    3416 => "000000000000000000",
    3417 => "000000000000000000",
    3418 => "000000000000000000",
    3419 => "000000000000000000",
    3420 => "000000000000000000",
    3421 => "000000000000000000",
    3422 => "000000000000000000",
    3423 => "000000000000000000",
    3424 => "000000000000000000",
    3425 => "000000000000000000",
    3426 => "000000000000000000",
    3427 => "000000000000000000",
    3428 => "000000000000000000",
    3429 => "000000000000000000",
    3430 => "000000000000000000",
    3431 => "000000000000000000",
    3432 => "000000000000000000",
    3433 => "000000000000000000",
    3434 => "000000000000000000",
    3435 => "000000000000000000",
    3436 => "000000000000000000",
    3437 => "000000000000000000",
    3438 => "000000000000000000",
    3439 => "000000000000000000",
    3440 => "000000000000000000",
    3441 => "000000000000000000",
    3442 => "000000000000000000",
    3443 => "000000000000000000",
    3444 => "000000000000000000",
    3445 => "000000000000000000",
    3446 => "000000000000000000",
    3447 => "000000000000000000",
    3448 => "000000000000000000",
    3449 => "000000000000000000",
    3450 => "000000000000000000",
    3451 => "000000000000000000",
    3452 => "000000000000000000",
    3453 => "000000000000000000",
    3454 => "000000000000000000",
    3455 => "000000000000000000",
    3456 => "000000000000000000",
    3457 => "000000000000000000",
    3458 => "000000000000000000",
    3459 => "000000000000000000",
    3460 => "000000000000000000",
    3461 => "000000000000000000",
    3462 => "000000000000000000",
    3463 => "000000000000000000",
    3464 => "000000000000000000",
    3465 => "000000000000000000",
    3466 => "000000000000000000",
    3467 => "000000000000000000",
    3468 => "000000000000000000",
    3469 => "000000000000000000",
    3470 => "000000000000000000",
    3471 => "000000000000000000",
    3472 => "000000000000000000",
    3473 => "000000000000000000",
    3474 => "000000000000000000",
    3475 => "000000000000000000",
    3476 => "000000000000000000",
    3477 => "000000000000000000",
    3478 => "000000000000000000",
    3479 => "000000000000000000",
    3480 => "000000000000000000",
    3481 => "000000000000000000",
    3482 => "000000000000000000",
    3483 => "000000000000000000",
    3484 => "000000000000000000",
    3485 => "000000000000000000",
    3486 => "000000000000000000",
    3487 => "000000000000000000",
    3488 => "000000000000000000",
    3489 => "000000000000000000",
    3490 => "000000000000000000",
    3491 => "000000000000000000",
    3492 => "000000000000000000",
    3493 => "000000000000000000",
    3494 => "000000000000000000",
    3495 => "000000000000000000",
    3496 => "000000000000000000",
    3497 => "000000000000000000",
    3498 => "000000000000000000",
    3499 => "000000000000000000",
    3500 => "000000000000000000",
    3501 => "000000000000000000",
    3502 => "000000000000000000",
    3503 => "000000000000000000",
    3504 => "000000000000000000",
    3505 => "000000000000000000",
    3506 => "000000000000000000",
    3507 => "000000000000000000",
    3508 => "000000000000000000",
    3509 => "000000000000000000",
    3510 => "000000000000000000",
    3511 => "000000000000000000",
    3512 => "000000000000000000",
    3513 => "000000000000000000",
    3514 => "000000000000000000",
    3515 => "000000000000000000",
    3516 => "000000000000000000",
    3517 => "000000000000000000",
    3518 => "000000000000000000",
    3519 => "000000000000000000",
    3520 => "000000000000000000",
    3521 => "000000000000000000",
    3522 => "000000000000000000",
    3523 => "000000000000000000",
    3524 => "000000000000000000",
    3525 => "000000000000000000",
    3526 => "000000000000000000",
    3527 => "000000000000000000",
    3528 => "000000000000000000",
    3529 => "000000000000000000",
    3530 => "000000000000000000",
    3531 => "000000000000000000",
    3532 => "000000000000000000",
    3533 => "000000000000000000",
    3534 => "000000000000000000",
    3535 => "000000000000000000",
    3536 => "000000000000000000",
    3537 => "000000000000000000",
    3538 => "000000000000000000",
    3539 => "000000000000000000",
    3540 => "000000000000000000",
    3541 => "000000000000000000",
    3542 => "000000000000000000",
    3543 => "000000000000000000",
    3544 => "000000000000000000",
    3545 => "000000000000000000",
    3546 => "000000000000000000",
    3547 => "000000000000000000",
    3548 => "000000000000000000",
    3549 => "000000000000000000",
    3550 => "000000000000000000",
    3551 => "000000000000000000",
    3552 => "000000000000000000",
    3553 => "000000000000000000",
    3554 => "000000000000000000",
    3555 => "000000000000000000",
    3556 => "000000000000000000",
    3557 => "000000000000000000",
    3558 => "000000000000000000",
    3559 => "000000000000000000",
    3560 => "000000000000000000",
    3561 => "000000000000000000",
    3562 => "000000000000000000",
    3563 => "000000000000000000",
    3564 => "000000000000000000",
    3565 => "000000000000000000",
    3566 => "000000000000000000",
    3567 => "000000000000000000",
    3568 => "000000000000000000",
    3569 => "000000000000000000",
    3570 => "000000000000000000",
    3571 => "000000000000000000",
    3572 => "000000000000000000",
    3573 => "000000000000000000",
    3574 => "000000000000000000",
    3575 => "000000000000000000",
    3576 => "000000000000000000",
    3577 => "000000000000000000",
    3578 => "000000000000000000",
    3579 => "000000000000000000",
    3580 => "000000000000000000",
    3581 => "000000000000000000",
    3582 => "000000000000000000",
    3583 => "000000000000000000",
    3584 => "000000000000000000",
    3585 => "000000000000000000",
    3586 => "000000000000000000",
    3587 => "000000000000000000",
    3588 => "000000000000000000",
    3589 => "000000000000000000",
    3590 => "000000000000000000",
    3591 => "000000000000000000",
    3592 => "000000000000000000",
    3593 => "000000000000000000",
    3594 => "000000000000000000",
    3595 => "000000000000000000",
    3596 => "000000000000000000",
    3597 => "000000000000000000",
    3598 => "000000000000000000",
    3599 => "000000000000000000",
    3600 => "000000000000000000",
    3601 => "000000000000000000",
    3602 => "000000000000000000",
    3603 => "000000000000000000",
    3604 => "000000000000000000",
    3605 => "000000000000000000",
    3606 => "000000000000000000",
    3607 => "000000000000000000",
    3608 => "000000000000000000",
    3609 => "000000000000000000",
    3610 => "000000000000000000",
    3611 => "000000000000000000",
    3612 => "000000000000000000",
    3613 => "000000000000000000",
    3614 => "000000000000000000",
    3615 => "000000000000000000",
    3616 => "000000000000000000",
    3617 => "000000000000000000",
    3618 => "000000000000000000",
    3619 => "000000000000000000",
    3620 => "000000000000000000",
    3621 => "000000000000000000",
    3622 => "000000000000000000",
    3623 => "000000000000000000",
    3624 => "000000000000000000",
    3625 => "000000000000000000",
    3626 => "000000000000000000",
    3627 => "000000000000000000",
    3628 => "000000000000000000",
    3629 => "000000000000000000",
    3630 => "000000000000000000",
    3631 => "000000000000000000",
    3632 => "000000000000000000",
    3633 => "000000000000000000",
    3634 => "000000000000000000",
    3635 => "000000000000000000",
    3636 => "000000000000000000",
    3637 => "000000000000000000",
    3638 => "000000000000000000",
    3639 => "000000000000000000",
    3640 => "000000000000000000",
    3641 => "000000000000000000",
    3642 => "000000000000000000",
    3643 => "000000000000000000",
    3644 => "000000000000000000",
    3645 => "000000000000000000",
    3646 => "000000000000000000",
    3647 => "000000000000000000",
    3648 => "000000000000000000",
    3649 => "000000000000000000",
    3650 => "000000000000000000",
    3651 => "000000000000000000",
    3652 => "000000000000000000",
    3653 => "000000000000000000",
    3654 => "000000000000000000",
    3655 => "000000000000000000",
    3656 => "000000000000000000",
    3657 => "000000000000000000",
    3658 => "000000000000000000",
    3659 => "000000000000000000",
    3660 => "000000000000000000",
    3661 => "000000000000000000",
    3662 => "000000000000000000",
    3663 => "000000000000000000",
    3664 => "000000000000000000",
    3665 => "000000000000000000",
    3666 => "000000000000000000",
    3667 => "000000000000000000",
    3668 => "000000000000000000",
    3669 => "000000000000000000",
    3670 => "000000000000000000",
    3671 => "000000000000000000",
    3672 => "000000000000000000",
    3673 => "000000000000000000",
    3674 => "000000000000000000",
    3675 => "000000000000000000",
    3676 => "000000000000000000",
    3677 => "000000000000000000",
    3678 => "000000000000000000",
    3679 => "000000000000000000",
    3680 => "000000000000000000",
    3681 => "000000000000000000",
    3682 => "000000000000000000",
    3683 => "000000000000000000",
    3684 => "000000000000000000",
    3685 => "000000000000000000",
    3686 => "000000000000000000",
    3687 => "000000000000000000",
    3688 => "000000000000000000",
    3689 => "000000000000000000",
    3690 => "000000000000000000",
    3691 => "000000000000000000",
    3692 => "000000000000000000",
    3693 => "000000000000000000",
    3694 => "000000000000000000",
    3695 => "000000000000000000",
    3696 => "000000000000000000",
    3697 => "000000000000000000",
    3698 => "000000000000000000",
    3699 => "000000000000000000",
    3700 => "000000000000000000",
    3701 => "000000000000000000",
    3702 => "000000000000000000",
    3703 => "000000000000000000",
    3704 => "000000000000000000",
    3705 => "000000000000000000",
    3706 => "000000000000000000",
    3707 => "000000000000000000",
    3708 => "000000000000000000",
    3709 => "000000000000000000",
    3710 => "000000000000000000",
    3711 => "000000000000000000",
    3712 => "000000000000000000",
    3713 => "000000000000000000",
    3714 => "000000000000000000",
    3715 => "000000000000000000",
    3716 => "000000000000000000",
    3717 => "000000000000000000",
    3718 => "000000000000000000",
    3719 => "000000000000000000",
    3720 => "000000000000000000",
    3721 => "000000000000000000",
    3722 => "000000000000000000",
    3723 => "000000000000000000",
    3724 => "000000000000000000",
    3725 => "000000000000000000",
    3726 => "000000000000000000",
    3727 => "000000000000000000",
    3728 => "000000000000000000",
    3729 => "000000000000000000",
    3730 => "000000000000000000",
    3731 => "000000000000000000",
    3732 => "000000000000000000",
    3733 => "000000000000000000",
    3734 => "000000000000000000",
    3735 => "000000000000000000",
    3736 => "000000000000000000",
    3737 => "000000000000000000",
    3738 => "000000000000000000",
    3739 => "000000000000000000",
    3740 => "000000000000000000",
    3741 => "000000000000000000",
    3742 => "000000000000000000",
    3743 => "000000000000000000",
    3744 => "000000000000000000",
    3745 => "000000000000000000",
    3746 => "000000000000000000",
    3747 => "000000000000000000",
    3748 => "000000000000000000",
    3749 => "000000000000000000",
    3750 => "000000000000000000",
    3751 => "000000000000000000",
    3752 => "000000000000000000",
    3753 => "000000000000000000",
    3754 => "000000000000000000",
    3755 => "000000000000000000",
    3756 => "000000000000000000",
    3757 => "000000000000000000",
    3758 => "000000000000000000",
    3759 => "000000000000000000",
    3760 => "000000000000000000",
    3761 => "000000000000000000",
    3762 => "000000000000000000",
    3763 => "000000000000000000",
    3764 => "000000000000000000",
    3765 => "000000000000000000",
    3766 => "000000000000000000",
    3767 => "000000000000000000",
    3768 => "000000000000000000",
    3769 => "000000000000000000",
    3770 => "000000000000000000",
    3771 => "000000000000000000",
    3772 => "000000000000000000",
    3773 => "000000000000000000",
    3774 => "000000000000000000",
    3775 => "000000000000000000",
    3776 => "000000000000000000",
    3777 => "000000000000000000",
    3778 => "000000000000000000",
    3779 => "000000000000000000",
    3780 => "000000000000000000",
    3781 => "000000000000000000",
    3782 => "000000000000000000",
    3783 => "000000000000000000",
    3784 => "000000000000000000",
    3785 => "000000000000000000",
    3786 => "000000000000000000",
    3787 => "000000000000000000",
    3788 => "000000000000000000",
    3789 => "000000000000000000",
    3790 => "000000000000000000",
    3791 => "000000000000000000",
    3792 => "000000000000000000",
    3793 => "000000000000000000",
    3794 => "000000000000000000",
    3795 => "000000000000000000",
    3796 => "000000000000000000",
    3797 => "000000000000000000",
    3798 => "000000000000000000",
    3799 => "000000000000000000",
    3800 => "000000000000000000",
    3801 => "000000000000000000",
    3802 => "000000000000000000",
    3803 => "000000000000000000",
    3804 => "000000000000000000",
    3805 => "000000000000000000",
    3806 => "000000000000000000",
    3807 => "000000000000000000",
    3808 => "000000000000000000",
    3809 => "000000000000000000",
    3810 => "000000000000000000",
    3811 => "000000000000000000",
    3812 => "000000000000000000",
    3813 => "000000000000000000",
    3814 => "000000000000000000",
    3815 => "000000000000000000",
    3816 => "000000000000000000",
    3817 => "000000000000000000",
    3818 => "000000000000000000",
    3819 => "000000000000000000",
    3820 => "000000000000000000",
    3821 => "000000000000000000",
    3822 => "000000000000000000",
    3823 => "000000000000000000",
    3824 => "000000000000000000",
    3825 => "000000000000000000",
    3826 => "000000000000000000",
    3827 => "000000000000000000",
    3828 => "000000000000000000",
    3829 => "000000000000000000",
    3830 => "000000000000000000",
    3831 => "000000000000000000",
    3832 => "000000000000000000",
    3833 => "000000000000000000",
    3834 => "000000000000000000",
    3835 => "000000000000000000",
    3836 => "000000000000000000",
    3837 => "000000000000000000",
    3838 => "000000000000000000",
    3839 => "000000000000000000",
    3840 => "000000000000000000",
    3841 => "000000000000000000",
    3842 => "000000000000000000",
    3843 => "000000000000000000",
    3844 => "000000000000000000",
    3845 => "000000000000000000",
    3846 => "000000000000000000",
    3847 => "000000000000000000",
    3848 => "000000000000000000",
    3849 => "000000000000000000",
    3850 => "000000000000000000",
    3851 => "000000000000000000",
    3852 => "000000000000000000",
    3853 => "000000000000000000",
    3854 => "000000000000000000",
    3855 => "000000000000000000",
    3856 => "000000000000000000",
    3857 => "000000000000000000",
    3858 => "000000000000000000",
    3859 => "000000000000000000",
    3860 => "000000000000000000",
    3861 => "000000000000000000",
    3862 => "000000000000000000",
    3863 => "000000000000000000",
    3864 => "000000000000000000",
    3865 => "000000000000000000",
    3866 => "000000000000000000",
    3867 => "000000000000000000",
    3868 => "000000000000000000",
    3869 => "000000000000000000",
    3870 => "000000000000000000",
    3871 => "000000000000000000",
    3872 => "000000000000000000",
    3873 => "000000000000000000",
    3874 => "000000000000000000",
    3875 => "000000000000000000",
    3876 => "000000000000000000",
    3877 => "000000000000000000",
    3878 => "000000000000000000",
    3879 => "000000000000000000",
    3880 => "000000000000000000",
    3881 => "000000000000000000",
    3882 => "000000000000000000",
    3883 => "000000000000000000",
    3884 => "000000000000000000",
    3885 => "000000000000000000",
    3886 => "000000000000000000",
    3887 => "000000000000000000",
    3888 => "000000000000000000",
    3889 => "000000000000000000",
    3890 => "000000000000000000",
    3891 => "000000000000000000",
    3892 => "000000000000000000",
    3893 => "000000000000000000",
    3894 => "000000000000000000",
    3895 => "000000000000000000",
    3896 => "000000000000000000",
    3897 => "000000000000000000",
    3898 => "000000000000000000",
    3899 => "000000000000000000",
    3900 => "000000000000000000",
    3901 => "000000000000000000",
    3902 => "000000000000000000",
    3903 => "000000000000000000",
    3904 => "000000000000000000",
    3905 => "000000000000000000",
    3906 => "000000000000000000",
    3907 => "000000000000000000",
    3908 => "000000000000000000",
    3909 => "000000000000000000",
    3910 => "000000000000000000",
    3911 => "000000000000000000",
    3912 => "000000000000000000",
    3913 => "000000000000000000",
    3914 => "000000000000000000",
    3915 => "000000000000000000",
    3916 => "000000000000000000",
    3917 => "000000000000000000",
    3918 => "000000000000000000",
    3919 => "000000000000000000",
    3920 => "000000000000000000",
    3921 => "000000000000000000",
    3922 => "000000000000000000",
    3923 => "000000000000000000",
    3924 => "000000000000000000",
    3925 => "000000000000000000",
    3926 => "000000000000000000",
    3927 => "000000000000000000",
    3928 => "000000000000000000",
    3929 => "000000000000000000",
    3930 => "000000000000000000",
    3931 => "000000000000000000",
    3932 => "000000000000000000",
    3933 => "000000000000000000",
    3934 => "000000000000000000",
    3935 => "000000000000000000",
    3936 => "000000000000000000",
    3937 => "000000000000000000",
    3938 => "000000000000000000",
    3939 => "000000000000000000",
    3940 => "000000000000000000",
    3941 => "000000000000000000",
    3942 => "000000000000000000",
    3943 => "000000000000000000",
    3944 => "000000000000000000",
    3945 => "000000000000000000",
    3946 => "000000000000000000",
    3947 => "000000000000000000",
    3948 => "000000000000000000",
    3949 => "000000000000000000",
    3950 => "000000000000000000",
    3951 => "000000000000000000",
    3952 => "000000000000000000",
    3953 => "000000000000000000",
    3954 => "000000000000000000",
    3955 => "000000000000000000",
    3956 => "000000000000000000",
    3957 => "000000000000000000",
    3958 => "000000000000000000",
    3959 => "000000000000000000",
    3960 => "000000000000000000",
    3961 => "000000000000000000",
    3962 => "000000000000000000",
    3963 => "000000000000000000",
    3964 => "000000000000000000",
    3965 => "000000000000000000",
    3966 => "000000000000000000",
    3967 => "000000000000000000",
    3968 => "000000000000000000",
    3969 => "000000000000000000",
    3970 => "000000000000000000",
    3971 => "000000000000000000",
    3972 => "000000000000000000",
    3973 => "000000000000000000",
    3974 => "000000000000000000",
    3975 => "000000000000000000",
    3976 => "000000000000000000",
    3977 => "000000000000000000",
    3978 => "000000000000000000",
    3979 => "000000000000000000",
    3980 => "000000000000000000",
    3981 => "000000000000000000",
    3982 => "000000000000000000",
    3983 => "000000000000000000",
    3984 => "000000000000000000",
    3985 => "000000000000000000",
    3986 => "000000000000000000",
    3987 => "000000000000000000",
    3988 => "000000000000000000",
    3989 => "000000000000000000",
    3990 => "000000000000000000",
    3991 => "000000000000000000",
    3992 => "000000000000000000",
    3993 => "000000000000000000",
    3994 => "000000000000000000",
    3995 => "000000000000000000",
    3996 => "000000000000000000",
    3997 => "000000000000000000",
    3998 => "000000000000000000",
    3999 => "000000000000000000",
    4000 => "000000000000000000",
    4001 => "000000000000000000",
    4002 => "000000000000000000",
    4003 => "000000000000000000",
    4004 => "000000000000000000",
    4005 => "000000000000000000",
    4006 => "000000000000000000",
    4007 => "000000000000000000",
    4008 => "000000000000000000",
    4009 => "000000000000000000",
    4010 => "000000000000000000",
    4011 => "000000000000000000",
    4012 => "000000000000000000",
    4013 => "000000000000000000",
    4014 => "000000000000000000",
    4015 => "000000000000000000",
    4016 => "000000000000000000",
    4017 => "000000000000000000",
    4018 => "000000000000000000",
    4019 => "000000000000000000",
    4020 => "000000000000000000",
    4021 => "000000000000000000",
    4022 => "000000000000000000",
    4023 => "000000000000000000",
    4024 => "000000000000000000",
    4025 => "000000000000000000",
    4026 => "000000000000000000",
    4027 => "000000000000000000",
    4028 => "000000000000000000",
    4029 => "000000000000000000",
    4030 => "000000000000000000",
    4031 => "000000000000000000",
    4032 => "000000000000000000",
    4033 => "000000000000000000",
    4034 => "000000000000000000",
    4035 => "000000000000000000",
    4036 => "000000000000000000",
    4037 => "000000000000000000",
    4038 => "000000000000000000",
    4039 => "000000000000000000",
    4040 => "000000000000000000",
    4041 => "000000000000000000",
    4042 => "000000000000000000",
    4043 => "000000000000000000",
    4044 => "000000000000000000",
    4045 => "000000000000000000",
    4046 => "000000000000000000",
    4047 => "000000000000000000",
    4048 => "000000000000000000",
    4049 => "000000000000000000",
    4050 => "000000000000000000",
    4051 => "000000000000000000",
    4052 => "000000000000000000",
    4053 => "000000000000000000",
    4054 => "000000000000000000",
    4055 => "000000000000000000",
    4056 => "000000000000000000",
    4057 => "000000000000000000",
    4058 => "000000000000000000",
    4059 => "000000000000000000",
    4060 => "000000000000000000",
    4061 => "000000000000000000",
    4062 => "000000000000000000",
    4063 => "000000000000000000",
    4064 => "000000000000000000",
    4065 => "000000000000000000",
    4066 => "000000000000000000",
    4067 => "000000000000000000",
    4068 => "000000000000000000",
    4069 => "000000000000000000",
    4070 => "000000000000000000",
    4071 => "000000000000000000",
    4072 => "000000000000000000",
    4073 => "000000000000000000",
    4074 => "000000000000000000",
    4075 => "000000000000000000",
    4076 => "000000000000000000",
    4077 => "000000000000000000",
    4078 => "000000000000000000",
    4079 => "000000000000000000",
    4080 => "000000000000000000",
    4081 => "000000000000000000",
    4082 => "000000000000000000",
    4083 => "000000000000000000",
    4084 => "000000000000000000",
    4085 => "000000000000000000",
    4086 => "000000000000000000",
    4087 => "000000000000000000",
    4088 => "000000000000000000",
    4089 => "000000000000000000",
    4090 => "000000000000000000",
    4091 => "000000000000000000",
    4092 => "000000000000000000",
    4093 => "000000000000000000",
    4094 => "000000000000000000",
    4095 => "000000000000000000" );
end package gasm_text;
